
module testrom (i_clock, i_cs, i_addr, o_data);
	input wire i_clock;
	input wire i_cs;
	input wire[14:0] i_addr;
	output wire[7:0] o_data = i_cs ? data : {8{1'bZ}};
	
	reg[7:0] data;
	
	always @(posedge i_clock) 
	begin
		case(i_addr)
			15'h00000000 : data <= 8'b10101001 ;
			15'h00000001 : data <= 8'b01001000 ;
			15'h00000002 : data <= 8'b10001101 ;
			15'h00000003 : data <= 8'b00000000 ;
			15'h00000004 : data <= 8'b01111110 ;
			15'h00000005 : data <= 8'b10101001 ;
			15'h00000006 : data <= 8'b01100101 ;
			15'h00000007 : data <= 8'b10001101 ;
			15'h00000008 : data <= 8'b00000001 ;
			15'h00000009 : data <= 8'b01111110 ;
			15'h0000000A : data <= 8'b10101001 ;
			15'h0000000B : data <= 8'b01101100 ;
			15'h0000000C : data <= 8'b10001101 ;
			15'h0000000D : data <= 8'b00000010 ;
			15'h0000000E : data <= 8'b01111110 ;
			15'h0000000F : data <= 8'b10101001 ;
			15'h00000010 : data <= 8'b01101100 ;
			15'h00000011 : data <= 8'b10001101 ;
			15'h00000012 : data <= 8'b00000011 ;
			15'h00000013 : data <= 8'b01111110 ;
			15'h00000014 : data <= 8'b10101001 ;
			15'h00000015 : data <= 8'b01101111 ;
			15'h00000016 : data <= 8'b10001101 ;
			15'h00000017 : data <= 8'b00000100 ;
			15'h00000018 : data <= 8'b01111110 ;
			15'h00000019 : data <= 8'b10101001 ;
			15'h0000001A : data <= 8'b00100000 ;
			15'h0000001B : data <= 8'b10001101 ;
			15'h0000001C : data <= 8'b00000101 ;
			15'h0000001D : data <= 8'b01111110 ;
			15'h0000001E : data <= 8'b10101001 ;
			15'h0000001F : data <= 8'b01010111 ;
			15'h00000020 : data <= 8'b10001101 ;
			15'h00000021 : data <= 8'b00000110 ;
			15'h00000022 : data <= 8'b01111110 ;
			15'h00000023 : data <= 8'b10101001 ;
			15'h00000024 : data <= 8'b01101111 ;
			15'h00000025 : data <= 8'b10001101 ;
			15'h00000026 : data <= 8'b00000111 ;
			15'h00000027 : data <= 8'b01111110 ;
			15'h00000028 : data <= 8'b10101001 ;
			15'h00000029 : data <= 8'b01110010 ;
			15'h0000002A : data <= 8'b10001101 ;
			15'h0000002B : data <= 8'b00001000 ;
			15'h0000002C : data <= 8'b01111110 ;
			15'h0000002D : data <= 8'b10101001 ;
			15'h0000002E : data <= 8'b01101100 ;
			15'h0000002F : data <= 8'b10001101 ;
			15'h00000030 : data <= 8'b00001001 ;
			15'h00000031 : data <= 8'b01111110 ;
			15'h00000032 : data <= 8'b10101001 ;
			15'h00000033 : data <= 8'b01100100 ;
			15'h00000034 : data <= 8'b10001101 ;
			15'h00000035 : data <= 8'b00001010 ;
			15'h00000036 : data <= 8'b01111110 ;
			15'h00000037 : data <= 8'b10101001 ;
			15'h00000038 : data <= 8'b00100001 ;
			15'h00000039 : data <= 8'b10001101 ;
			15'h0000003A : data <= 8'b00001011 ;
			15'h0000003B : data <= 8'b01111110 ;
			15'h0000003C : data <= 8'b11110010 ;
			15'h0000003D : data <= 8'b00000000 ;
			15'h0000003E : data <= 8'b00000000 ;
			15'h0000003F : data <= 8'b00000000 ;
			15'h00000040 : data <= 8'b00000000 ;
			15'h00000041 : data <= 8'b00000000 ;
			15'h00000042 : data <= 8'b00000000 ;
			15'h00000043 : data <= 8'b00000000 ;
			15'h00000044 : data <= 8'b00000000 ;
			15'h00000045 : data <= 8'b00000000 ;
			15'h00000046 : data <= 8'b00000000 ;
			15'h00000047 : data <= 8'b00000000 ;
			15'h00000048 : data <= 8'b00000000 ;
			15'h00000049 : data <= 8'b00000000 ;
			15'h0000004A : data <= 8'b00000000 ;
			15'h0000004B : data <= 8'b00000000 ;
			15'h0000004C : data <= 8'b00000000 ;
			15'h0000004D : data <= 8'b00000000 ;
			15'h0000004E : data <= 8'b00000000 ;
			15'h0000004F : data <= 8'b00000000 ;
			15'h00000050 : data <= 8'b00000000 ;
			15'h00000051 : data <= 8'b00000000 ;
			15'h00000052 : data <= 8'b00000000 ;
			15'h00000053 : data <= 8'b00000000 ;
			15'h00000054 : data <= 8'b00000000 ;
			15'h00000055 : data <= 8'b00000000 ;
			15'h00000056 : data <= 8'b00000000 ;
			15'h00000057 : data <= 8'b00000000 ;
			15'h00000058 : data <= 8'b00000000 ;
			15'h00000059 : data <= 8'b00000000 ;
			15'h0000005A : data <= 8'b00000000 ;
			15'h0000005B : data <= 8'b00000000 ;
			15'h0000005C : data <= 8'b00000000 ;
			15'h0000005D : data <= 8'b00000000 ;
			15'h0000005E : data <= 8'b00000000 ;
			15'h0000005F : data <= 8'b00000000 ;
			15'h00000060 : data <= 8'b00000000 ;
			15'h00000061 : data <= 8'b00000000 ;
			15'h00000062 : data <= 8'b00000000 ;
			15'h00000063 : data <= 8'b00000000 ;
			15'h00000064 : data <= 8'b00000000 ;
			15'h00000065 : data <= 8'b00000000 ;
			15'h00000066 : data <= 8'b00000000 ;
			15'h00000067 : data <= 8'b00000000 ;
			15'h00000068 : data <= 8'b00000000 ;
			15'h00000069 : data <= 8'b00000000 ;
			15'h0000006A : data <= 8'b00000000 ;
			15'h0000006B : data <= 8'b00000000 ;
			15'h0000006C : data <= 8'b00000000 ;
			15'h0000006D : data <= 8'b00000000 ;
			15'h0000006E : data <= 8'b00000000 ;
			15'h0000006F : data <= 8'b00000000 ;
			15'h00000070 : data <= 8'b00000000 ;
			15'h00000071 : data <= 8'b00000000 ;
			15'h00000072 : data <= 8'b00000000 ;
			15'h00000073 : data <= 8'b00000000 ;
			15'h00000074 : data <= 8'b00000000 ;
			15'h00000075 : data <= 8'b00000000 ;
			15'h00000076 : data <= 8'b00000000 ;
			15'h00000077 : data <= 8'b00000000 ;
			15'h00000078 : data <= 8'b00000000 ;
			15'h00000079 : data <= 8'b00000000 ;
			15'h0000007A : data <= 8'b00000000 ;
			15'h0000007B : data <= 8'b00000000 ;
			15'h0000007C : data <= 8'b00000000 ;
			15'h0000007D : data <= 8'b00000000 ;
			15'h0000007E : data <= 8'b00000000 ;
			15'h0000007F : data <= 8'b00000000 ;
			15'h00000080 : data <= 8'b00000000 ;
			15'h00000081 : data <= 8'b00000000 ;
			15'h00000082 : data <= 8'b00000000 ;
			15'h00000083 : data <= 8'b00000000 ;
			15'h00000084 : data <= 8'b00000000 ;
			15'h00000085 : data <= 8'b00000000 ;
			15'h00000086 : data <= 8'b00000000 ;
			15'h00000087 : data <= 8'b00000000 ;
			15'h00000088 : data <= 8'b00000000 ;
			15'h00000089 : data <= 8'b00000000 ;
			15'h0000008A : data <= 8'b00000000 ;
			15'h0000008B : data <= 8'b00000000 ;
			15'h0000008C : data <= 8'b00000000 ;
			15'h0000008D : data <= 8'b00000000 ;
			15'h0000008E : data <= 8'b00000000 ;
			15'h0000008F : data <= 8'b00000000 ;
			15'h00000090 : data <= 8'b00000000 ;
			15'h00000091 : data <= 8'b00000000 ;
			15'h00000092 : data <= 8'b00000000 ;
			15'h00000093 : data <= 8'b00000000 ;
			15'h00000094 : data <= 8'b00000000 ;
			15'h00000095 : data <= 8'b00000000 ;
			15'h00000096 : data <= 8'b00000000 ;
			15'h00000097 : data <= 8'b00000000 ;
			15'h00000098 : data <= 8'b00000000 ;
			15'h00000099 : data <= 8'b00000000 ;
			15'h0000009A : data <= 8'b00000000 ;
			15'h0000009B : data <= 8'b00000000 ;
			15'h0000009C : data <= 8'b00000000 ;
			15'h0000009D : data <= 8'b00000000 ;
			15'h0000009E : data <= 8'b00000000 ;
			15'h0000009F : data <= 8'b00000000 ;
			15'h000000A0 : data <= 8'b00000000 ;
			15'h000000A1 : data <= 8'b00000000 ;
			15'h000000A2 : data <= 8'b00000000 ;
			15'h000000A3 : data <= 8'b00000000 ;
			15'h000000A4 : data <= 8'b00000000 ;
			15'h000000A5 : data <= 8'b00000000 ;
			15'h000000A6 : data <= 8'b00000000 ;
			15'h000000A7 : data <= 8'b00000000 ;
			15'h000000A8 : data <= 8'b00000000 ;
			15'h000000A9 : data <= 8'b00000000 ;
			15'h000000AA : data <= 8'b00000000 ;
			15'h000000AB : data <= 8'b00000000 ;
			15'h000000AC : data <= 8'b00000000 ;
			15'h000000AD : data <= 8'b00000000 ;
			15'h000000AE : data <= 8'b00000000 ;
			15'h000000AF : data <= 8'b00000000 ;
			15'h000000B0 : data <= 8'b00000000 ;
			15'h000000B1 : data <= 8'b00000000 ;
			15'h000000B2 : data <= 8'b00000000 ;
			15'h000000B3 : data <= 8'b00000000 ;
			15'h000000B4 : data <= 8'b00000000 ;
			15'h000000B5 : data <= 8'b00000000 ;
			15'h000000B6 : data <= 8'b00000000 ;
			15'h000000B7 : data <= 8'b00000000 ;
			15'h000000B8 : data <= 8'b00000000 ;
			15'h000000B9 : data <= 8'b00000000 ;
			15'h000000BA : data <= 8'b00000000 ;
			15'h000000BB : data <= 8'b00000000 ;
			15'h000000BC : data <= 8'b00000000 ;
			15'h000000BD : data <= 8'b00000000 ;
			15'h000000BE : data <= 8'b00000000 ;
			15'h000000BF : data <= 8'b00000000 ;
			15'h000000C0 : data <= 8'b00000000 ;
			15'h000000C1 : data <= 8'b00000000 ;
			15'h000000C2 : data <= 8'b00000000 ;
			15'h000000C3 : data <= 8'b00000000 ;
			15'h000000C4 : data <= 8'b00000000 ;
			15'h000000C5 : data <= 8'b00000000 ;
			15'h000000C6 : data <= 8'b00000000 ;
			15'h000000C7 : data <= 8'b00000000 ;
			15'h000000C8 : data <= 8'b00000000 ;
			15'h000000C9 : data <= 8'b00000000 ;
			15'h000000CA : data <= 8'b00000000 ;
			15'h000000CB : data <= 8'b00000000 ;
			15'h000000CC : data <= 8'b00000000 ;
			15'h000000CD : data <= 8'b00000000 ;
			15'h000000CE : data <= 8'b00000000 ;
			15'h000000CF : data <= 8'b00000000 ;
			15'h000000D0 : data <= 8'b00000000 ;
			15'h000000D1 : data <= 8'b00000000 ;
			15'h000000D2 : data <= 8'b00000000 ;
			15'h000000D3 : data <= 8'b00000000 ;
			15'h000000D4 : data <= 8'b00000000 ;
			15'h000000D5 : data <= 8'b00000000 ;
			15'h000000D6 : data <= 8'b00000000 ;
			15'h000000D7 : data <= 8'b00000000 ;
			15'h000000D8 : data <= 8'b00000000 ;
			15'h000000D9 : data <= 8'b00000000 ;
			15'h000000DA : data <= 8'b00000000 ;
			15'h000000DB : data <= 8'b00000000 ;
			15'h000000DC : data <= 8'b00000000 ;
			15'h000000DD : data <= 8'b00000000 ;
			15'h000000DE : data <= 8'b00000000 ;
			15'h000000DF : data <= 8'b00000000 ;
			15'h000000E0 : data <= 8'b00000000 ;
			15'h000000E1 : data <= 8'b00000000 ;
			15'h000000E2 : data <= 8'b00000000 ;
			15'h000000E3 : data <= 8'b00000000 ;
			15'h000000E4 : data <= 8'b00000000 ;
			15'h000000E5 : data <= 8'b00000000 ;
			15'h000000E6 : data <= 8'b00000000 ;
			15'h000000E7 : data <= 8'b00000000 ;
			15'h000000E8 : data <= 8'b00000000 ;
			15'h000000E9 : data <= 8'b00000000 ;
			15'h000000EA : data <= 8'b00000000 ;
			15'h000000EB : data <= 8'b00000000 ;
			15'h000000EC : data <= 8'b00000000 ;
			15'h000000ED : data <= 8'b00000000 ;
			15'h000000EE : data <= 8'b00000000 ;
			15'h000000EF : data <= 8'b00000000 ;
			15'h000000F0 : data <= 8'b00000000 ;
			15'h000000F1 : data <= 8'b00000000 ;
			15'h000000F2 : data <= 8'b00000000 ;
			15'h000000F3 : data <= 8'b00000000 ;
			15'h000000F4 : data <= 8'b00000000 ;
			15'h000000F5 : data <= 8'b00000000 ;
			15'h000000F6 : data <= 8'b00000000 ;
			15'h000000F7 : data <= 8'b00000000 ;
			15'h000000F8 : data <= 8'b00000000 ;
			15'h000000F9 : data <= 8'b00000000 ;
			15'h000000FA : data <= 8'b00000000 ;
			15'h000000FB : data <= 8'b00000000 ;
			15'h000000FC : data <= 8'b00000000 ;
			15'h000000FD : data <= 8'b00000000 ;
			15'h000000FE : data <= 8'b00000000 ;
			15'h000000FF : data <= 8'b00000000 ;
			15'h00000100 : data <= 8'b00000000 ;
			15'h00000101 : data <= 8'b00000000 ;
			15'h00000102 : data <= 8'b00000000 ;
			15'h00000103 : data <= 8'b00000000 ;
			15'h00000104 : data <= 8'b00000000 ;
			15'h00000105 : data <= 8'b00000000 ;
			15'h00000106 : data <= 8'b00000000 ;
			15'h00000107 : data <= 8'b00000000 ;
			15'h00000108 : data <= 8'b00000000 ;
			15'h00000109 : data <= 8'b00000000 ;
			15'h0000010A : data <= 8'b00000000 ;
			15'h0000010B : data <= 8'b00000000 ;
			15'h0000010C : data <= 8'b00000000 ;
			15'h0000010D : data <= 8'b00000000 ;
			15'h0000010E : data <= 8'b00000000 ;
			15'h0000010F : data <= 8'b00000000 ;
			15'h00000110 : data <= 8'b00000000 ;
			15'h00000111 : data <= 8'b00000000 ;
			15'h00000112 : data <= 8'b00000000 ;
			15'h00000113 : data <= 8'b00000000 ;
			15'h00000114 : data <= 8'b00000000 ;
			15'h00000115 : data <= 8'b00000000 ;
			15'h00000116 : data <= 8'b00000000 ;
			15'h00000117 : data <= 8'b00000000 ;
			15'h00000118 : data <= 8'b00000000 ;
			15'h00000119 : data <= 8'b00000000 ;
			15'h0000011A : data <= 8'b00000000 ;
			15'h0000011B : data <= 8'b00000000 ;
			15'h0000011C : data <= 8'b00000000 ;
			15'h0000011D : data <= 8'b00000000 ;
			15'h0000011E : data <= 8'b00000000 ;
			15'h0000011F : data <= 8'b00000000 ;
			15'h00000120 : data <= 8'b00000000 ;
			15'h00000121 : data <= 8'b00000000 ;
			15'h00000122 : data <= 8'b00000000 ;
			15'h00000123 : data <= 8'b00000000 ;
			15'h00000124 : data <= 8'b00000000 ;
			15'h00000125 : data <= 8'b00000000 ;
			15'h00000126 : data <= 8'b00000000 ;
			15'h00000127 : data <= 8'b00000000 ;
			15'h00000128 : data <= 8'b00000000 ;
			15'h00000129 : data <= 8'b00000000 ;
			15'h0000012A : data <= 8'b00000000 ;
			15'h0000012B : data <= 8'b00000000 ;
			15'h0000012C : data <= 8'b00000000 ;
			15'h0000012D : data <= 8'b00000000 ;
			15'h0000012E : data <= 8'b00000000 ;
			15'h0000012F : data <= 8'b00000000 ;
			15'h00000130 : data <= 8'b00000000 ;
			15'h00000131 : data <= 8'b00000000 ;
			15'h00000132 : data <= 8'b00000000 ;
			15'h00000133 : data <= 8'b00000000 ;
			15'h00000134 : data <= 8'b00000000 ;
			15'h00000135 : data <= 8'b00000000 ;
			15'h00000136 : data <= 8'b00000000 ;
			15'h00000137 : data <= 8'b00000000 ;
			15'h00000138 : data <= 8'b00000000 ;
			15'h00000139 : data <= 8'b00000000 ;
			15'h0000013A : data <= 8'b00000000 ;
			15'h0000013B : data <= 8'b00000000 ;
			15'h0000013C : data <= 8'b00000000 ;
			15'h0000013D : data <= 8'b00000000 ;
			15'h0000013E : data <= 8'b00000000 ;
			15'h0000013F : data <= 8'b00000000 ;
			15'h00000140 : data <= 8'b00000000 ;
			15'h00000141 : data <= 8'b00000000 ;
			15'h00000142 : data <= 8'b00000000 ;
			15'h00000143 : data <= 8'b00000000 ;
			15'h00000144 : data <= 8'b00000000 ;
			15'h00000145 : data <= 8'b00000000 ;
			15'h00000146 : data <= 8'b00000000 ;
			15'h00000147 : data <= 8'b00000000 ;
			15'h00000148 : data <= 8'b00000000 ;
			15'h00000149 : data <= 8'b00000000 ;
			15'h0000014A : data <= 8'b00000000 ;
			15'h0000014B : data <= 8'b00000000 ;
			15'h0000014C : data <= 8'b00000000 ;
			15'h0000014D : data <= 8'b00000000 ;
			15'h0000014E : data <= 8'b00000000 ;
			15'h0000014F : data <= 8'b00000000 ;
			15'h00000150 : data <= 8'b00000000 ;
			15'h00000151 : data <= 8'b00000000 ;
			15'h00000152 : data <= 8'b00000000 ;
			15'h00000153 : data <= 8'b00000000 ;
			15'h00000154 : data <= 8'b00000000 ;
			15'h00000155 : data <= 8'b00000000 ;
			15'h00000156 : data <= 8'b00000000 ;
			15'h00000157 : data <= 8'b00000000 ;
			15'h00000158 : data <= 8'b00000000 ;
			15'h00000159 : data <= 8'b00000000 ;
			15'h0000015A : data <= 8'b00000000 ;
			15'h0000015B : data <= 8'b00000000 ;
			15'h0000015C : data <= 8'b00000000 ;
			15'h0000015D : data <= 8'b00000000 ;
			15'h0000015E : data <= 8'b00000000 ;
			15'h0000015F : data <= 8'b00000000 ;
			15'h00000160 : data <= 8'b00000000 ;
			15'h00000161 : data <= 8'b00000000 ;
			15'h00000162 : data <= 8'b00000000 ;
			15'h00000163 : data <= 8'b00000000 ;
			15'h00000164 : data <= 8'b00000000 ;
			15'h00000165 : data <= 8'b00000000 ;
			15'h00000166 : data <= 8'b00000000 ;
			15'h00000167 : data <= 8'b00000000 ;
			15'h00000168 : data <= 8'b00000000 ;
			15'h00000169 : data <= 8'b00000000 ;
			15'h0000016A : data <= 8'b00000000 ;
			15'h0000016B : data <= 8'b00000000 ;
			15'h0000016C : data <= 8'b00000000 ;
			15'h0000016D : data <= 8'b00000000 ;
			15'h0000016E : data <= 8'b00000000 ;
			15'h0000016F : data <= 8'b00000000 ;
			15'h00000170 : data <= 8'b00000000 ;
			15'h00000171 : data <= 8'b00000000 ;
			15'h00000172 : data <= 8'b00000000 ;
			15'h00000173 : data <= 8'b00000000 ;
			15'h00000174 : data <= 8'b00000000 ;
			15'h00000175 : data <= 8'b00000000 ;
			15'h00000176 : data <= 8'b00000000 ;
			15'h00000177 : data <= 8'b00000000 ;
			15'h00000178 : data <= 8'b00000000 ;
			15'h00000179 : data <= 8'b00000000 ;
			15'h0000017A : data <= 8'b00000000 ;
			15'h0000017B : data <= 8'b00000000 ;
			15'h0000017C : data <= 8'b00000000 ;
			15'h0000017D : data <= 8'b00000000 ;
			15'h0000017E : data <= 8'b00000000 ;
			15'h0000017F : data <= 8'b00000000 ;
			15'h00000180 : data <= 8'b00000000 ;
			15'h00000181 : data <= 8'b00000000 ;
			15'h00000182 : data <= 8'b00000000 ;
			15'h00000183 : data <= 8'b00000000 ;
			15'h00000184 : data <= 8'b00000000 ;
			15'h00000185 : data <= 8'b00000000 ;
			15'h00000186 : data <= 8'b00000000 ;
			15'h00000187 : data <= 8'b00000000 ;
			15'h00000188 : data <= 8'b00000000 ;
			15'h00000189 : data <= 8'b00000000 ;
			15'h0000018A : data <= 8'b00000000 ;
			15'h0000018B : data <= 8'b00000000 ;
			15'h0000018C : data <= 8'b00000000 ;
			15'h0000018D : data <= 8'b00000000 ;
			15'h0000018E : data <= 8'b00000000 ;
			15'h0000018F : data <= 8'b00000000 ;
			15'h00000190 : data <= 8'b00000000 ;
			15'h00000191 : data <= 8'b00000000 ;
			15'h00000192 : data <= 8'b00000000 ;
			15'h00000193 : data <= 8'b00000000 ;
			15'h00000194 : data <= 8'b00000000 ;
			15'h00000195 : data <= 8'b00000000 ;
			15'h00000196 : data <= 8'b00000000 ;
			15'h00000197 : data <= 8'b00000000 ;
			15'h00000198 : data <= 8'b00000000 ;
			15'h00000199 : data <= 8'b00000000 ;
			15'h0000019A : data <= 8'b00000000 ;
			15'h0000019B : data <= 8'b00000000 ;
			15'h0000019C : data <= 8'b00000000 ;
			15'h0000019D : data <= 8'b00000000 ;
			15'h0000019E : data <= 8'b00000000 ;
			15'h0000019F : data <= 8'b00000000 ;
			15'h000001A0 : data <= 8'b00000000 ;
			15'h000001A1 : data <= 8'b00000000 ;
			15'h000001A2 : data <= 8'b00000000 ;
			15'h000001A3 : data <= 8'b00000000 ;
			15'h000001A4 : data <= 8'b00000000 ;
			15'h000001A5 : data <= 8'b00000000 ;
			15'h000001A6 : data <= 8'b00000000 ;
			15'h000001A7 : data <= 8'b00000000 ;
			15'h000001A8 : data <= 8'b00000000 ;
			15'h000001A9 : data <= 8'b00000000 ;
			15'h000001AA : data <= 8'b00000000 ;
			15'h000001AB : data <= 8'b00000000 ;
			15'h000001AC : data <= 8'b00000000 ;
			15'h000001AD : data <= 8'b00000000 ;
			15'h000001AE : data <= 8'b00000000 ;
			15'h000001AF : data <= 8'b00000000 ;
			15'h000001B0 : data <= 8'b00000000 ;
			15'h000001B1 : data <= 8'b00000000 ;
			15'h000001B2 : data <= 8'b00000000 ;
			15'h000001B3 : data <= 8'b00000000 ;
			15'h000001B4 : data <= 8'b00000000 ;
			15'h000001B5 : data <= 8'b00000000 ;
			15'h000001B6 : data <= 8'b00000000 ;
			15'h000001B7 : data <= 8'b00000000 ;
			15'h000001B8 : data <= 8'b00000000 ;
			15'h000001B9 : data <= 8'b00000000 ;
			15'h000001BA : data <= 8'b00000000 ;
			15'h000001BB : data <= 8'b00000000 ;
			15'h000001BC : data <= 8'b00000000 ;
			15'h000001BD : data <= 8'b00000000 ;
			15'h000001BE : data <= 8'b00000000 ;
			15'h000001BF : data <= 8'b00000000 ;
			15'h000001C0 : data <= 8'b00000000 ;
			15'h000001C1 : data <= 8'b00000000 ;
			15'h000001C2 : data <= 8'b00000000 ;
			15'h000001C3 : data <= 8'b00000000 ;
			15'h000001C4 : data <= 8'b00000000 ;
			15'h000001C5 : data <= 8'b00000000 ;
			15'h000001C6 : data <= 8'b00000000 ;
			15'h000001C7 : data <= 8'b00000000 ;
			15'h000001C8 : data <= 8'b00000000 ;
			15'h000001C9 : data <= 8'b00000000 ;
			15'h000001CA : data <= 8'b00000000 ;
			15'h000001CB : data <= 8'b00000000 ;
			15'h000001CC : data <= 8'b00000000 ;
			15'h000001CD : data <= 8'b00000000 ;
			15'h000001CE : data <= 8'b00000000 ;
			15'h000001CF : data <= 8'b00000000 ;
			15'h000001D0 : data <= 8'b00000000 ;
			15'h000001D1 : data <= 8'b00000000 ;
			15'h000001D2 : data <= 8'b00000000 ;
			15'h000001D3 : data <= 8'b00000000 ;
			15'h000001D4 : data <= 8'b00000000 ;
			15'h000001D5 : data <= 8'b00000000 ;
			15'h000001D6 : data <= 8'b00000000 ;
			15'h000001D7 : data <= 8'b00000000 ;
			15'h000001D8 : data <= 8'b00000000 ;
			15'h000001D9 : data <= 8'b00000000 ;
			15'h000001DA : data <= 8'b00000000 ;
			15'h000001DB : data <= 8'b00000000 ;
			15'h000001DC : data <= 8'b00000000 ;
			15'h000001DD : data <= 8'b00000000 ;
			15'h000001DE : data <= 8'b00000000 ;
			15'h000001DF : data <= 8'b00000000 ;
			15'h000001E0 : data <= 8'b00000000 ;
			15'h000001E1 : data <= 8'b00000000 ;
			15'h000001E2 : data <= 8'b00000000 ;
			15'h000001E3 : data <= 8'b00000000 ;
			15'h000001E4 : data <= 8'b00000000 ;
			15'h000001E5 : data <= 8'b00000000 ;
			15'h000001E6 : data <= 8'b00000000 ;
			15'h000001E7 : data <= 8'b00000000 ;
			15'h000001E8 : data <= 8'b00000000 ;
			15'h000001E9 : data <= 8'b00000000 ;
			15'h000001EA : data <= 8'b00000000 ;
			15'h000001EB : data <= 8'b00000000 ;
			15'h000001EC : data <= 8'b00000000 ;
			15'h000001ED : data <= 8'b00000000 ;
			15'h000001EE : data <= 8'b00000000 ;
			15'h000001EF : data <= 8'b00000000 ;
			15'h000001F0 : data <= 8'b00000000 ;
			15'h000001F1 : data <= 8'b00000000 ;
			15'h000001F2 : data <= 8'b00000000 ;
			15'h000001F3 : data <= 8'b00000000 ;
			15'h000001F4 : data <= 8'b00000000 ;
			15'h000001F5 : data <= 8'b00000000 ;
			15'h000001F6 : data <= 8'b00000000 ;
			15'h000001F7 : data <= 8'b00000000 ;
			15'h000001F8 : data <= 8'b00000000 ;
			15'h000001F9 : data <= 8'b00000000 ;
			15'h000001FA : data <= 8'b00000000 ;
			15'h000001FB : data <= 8'b00000000 ;
			15'h000001FC : data <= 8'b00000000 ;
			15'h000001FD : data <= 8'b00000000 ;
			15'h000001FE : data <= 8'b00000000 ;
			15'h000001FF : data <= 8'b00000000 ;
			15'h00000200 : data <= 8'b00000000 ;
			15'h00000201 : data <= 8'b00000000 ;
			15'h00000202 : data <= 8'b00000000 ;
			15'h00000203 : data <= 8'b00000000 ;
			15'h00000204 : data <= 8'b00000000 ;
			15'h00000205 : data <= 8'b00000000 ;
			15'h00000206 : data <= 8'b00000000 ;
			15'h00000207 : data <= 8'b00000000 ;
			15'h00000208 : data <= 8'b00000000 ;
			15'h00000209 : data <= 8'b00000000 ;
			15'h0000020A : data <= 8'b00000000 ;
			15'h0000020B : data <= 8'b00000000 ;
			15'h0000020C : data <= 8'b00000000 ;
			15'h0000020D : data <= 8'b00000000 ;
			15'h0000020E : data <= 8'b00000000 ;
			15'h0000020F : data <= 8'b00000000 ;
			15'h00000210 : data <= 8'b00000000 ;
			15'h00000211 : data <= 8'b00000000 ;
			15'h00000212 : data <= 8'b00000000 ;
			15'h00000213 : data <= 8'b00000000 ;
			15'h00000214 : data <= 8'b00000000 ;
			15'h00000215 : data <= 8'b00000000 ;
			15'h00000216 : data <= 8'b00000000 ;
			15'h00000217 : data <= 8'b00000000 ;
			15'h00000218 : data <= 8'b00000000 ;
			15'h00000219 : data <= 8'b00000000 ;
			15'h0000021A : data <= 8'b00000000 ;
			15'h0000021B : data <= 8'b00000000 ;
			15'h0000021C : data <= 8'b00000000 ;
			15'h0000021D : data <= 8'b00000000 ;
			15'h0000021E : data <= 8'b00000000 ;
			15'h0000021F : data <= 8'b00000000 ;
			15'h00000220 : data <= 8'b00000000 ;
			15'h00000221 : data <= 8'b00000000 ;
			15'h00000222 : data <= 8'b00000000 ;
			15'h00000223 : data <= 8'b00000000 ;
			15'h00000224 : data <= 8'b00000000 ;
			15'h00000225 : data <= 8'b00000000 ;
			15'h00000226 : data <= 8'b00000000 ;
			15'h00000227 : data <= 8'b00000000 ;
			15'h00000228 : data <= 8'b00000000 ;
			15'h00000229 : data <= 8'b00000000 ;
			15'h0000022A : data <= 8'b00000000 ;
			15'h0000022B : data <= 8'b00000000 ;
			15'h0000022C : data <= 8'b00000000 ;
			15'h0000022D : data <= 8'b00000000 ;
			15'h0000022E : data <= 8'b00000000 ;
			15'h0000022F : data <= 8'b00000000 ;
			15'h00000230 : data <= 8'b00000000 ;
			15'h00000231 : data <= 8'b00000000 ;
			15'h00000232 : data <= 8'b00000000 ;
			15'h00000233 : data <= 8'b00000000 ;
			15'h00000234 : data <= 8'b00000000 ;
			15'h00000235 : data <= 8'b00000000 ;
			15'h00000236 : data <= 8'b00000000 ;
			15'h00000237 : data <= 8'b00000000 ;
			15'h00000238 : data <= 8'b00000000 ;
			15'h00000239 : data <= 8'b00000000 ;
			15'h0000023A : data <= 8'b00000000 ;
			15'h0000023B : data <= 8'b00000000 ;
			15'h0000023C : data <= 8'b00000000 ;
			15'h0000023D : data <= 8'b00000000 ;
			15'h0000023E : data <= 8'b00000000 ;
			15'h0000023F : data <= 8'b00000000 ;
			15'h00000240 : data <= 8'b00000000 ;
			15'h00000241 : data <= 8'b00000000 ;
			15'h00000242 : data <= 8'b00000000 ;
			15'h00000243 : data <= 8'b00000000 ;
			15'h00000244 : data <= 8'b00000000 ;
			15'h00000245 : data <= 8'b00000000 ;
			15'h00000246 : data <= 8'b00000000 ;
			15'h00000247 : data <= 8'b00000000 ;
			15'h00000248 : data <= 8'b00000000 ;
			15'h00000249 : data <= 8'b00000000 ;
			15'h0000024A : data <= 8'b00000000 ;
			15'h0000024B : data <= 8'b00000000 ;
			15'h0000024C : data <= 8'b00000000 ;
			15'h0000024D : data <= 8'b00000000 ;
			15'h0000024E : data <= 8'b00000000 ;
			15'h0000024F : data <= 8'b00000000 ;
			15'h00000250 : data <= 8'b00000000 ;
			15'h00000251 : data <= 8'b00000000 ;
			15'h00000252 : data <= 8'b00000000 ;
			15'h00000253 : data <= 8'b00000000 ;
			15'h00000254 : data <= 8'b00000000 ;
			15'h00000255 : data <= 8'b00000000 ;
			15'h00000256 : data <= 8'b00000000 ;
			15'h00000257 : data <= 8'b00000000 ;
			15'h00000258 : data <= 8'b00000000 ;
			15'h00000259 : data <= 8'b00000000 ;
			15'h0000025A : data <= 8'b00000000 ;
			15'h0000025B : data <= 8'b00000000 ;
			15'h0000025C : data <= 8'b00000000 ;
			15'h0000025D : data <= 8'b00000000 ;
			15'h0000025E : data <= 8'b00000000 ;
			15'h0000025F : data <= 8'b00000000 ;
			15'h00000260 : data <= 8'b00000000 ;
			15'h00000261 : data <= 8'b00000000 ;
			15'h00000262 : data <= 8'b00000000 ;
			15'h00000263 : data <= 8'b00000000 ;
			15'h00000264 : data <= 8'b00000000 ;
			15'h00000265 : data <= 8'b00000000 ;
			15'h00000266 : data <= 8'b00000000 ;
			15'h00000267 : data <= 8'b00000000 ;
			15'h00000268 : data <= 8'b00000000 ;
			15'h00000269 : data <= 8'b00000000 ;
			15'h0000026A : data <= 8'b00000000 ;
			15'h0000026B : data <= 8'b00000000 ;
			15'h0000026C : data <= 8'b00000000 ;
			15'h0000026D : data <= 8'b00000000 ;
			15'h0000026E : data <= 8'b00000000 ;
			15'h0000026F : data <= 8'b00000000 ;
			15'h00000270 : data <= 8'b00000000 ;
			15'h00000271 : data <= 8'b00000000 ;
			15'h00000272 : data <= 8'b00000000 ;
			15'h00000273 : data <= 8'b00000000 ;
			15'h00000274 : data <= 8'b00000000 ;
			15'h00000275 : data <= 8'b00000000 ;
			15'h00000276 : data <= 8'b00000000 ;
			15'h00000277 : data <= 8'b00000000 ;
			15'h00000278 : data <= 8'b00000000 ;
			15'h00000279 : data <= 8'b00000000 ;
			15'h0000027A : data <= 8'b00000000 ;
			15'h0000027B : data <= 8'b00000000 ;
			15'h0000027C : data <= 8'b00000000 ;
			15'h0000027D : data <= 8'b00000000 ;
			15'h0000027E : data <= 8'b00000000 ;
			15'h0000027F : data <= 8'b00000000 ;
			15'h00000280 : data <= 8'b00000000 ;
			15'h00000281 : data <= 8'b00000000 ;
			15'h00000282 : data <= 8'b00000000 ;
			15'h00000283 : data <= 8'b00000000 ;
			15'h00000284 : data <= 8'b00000000 ;
			15'h00000285 : data <= 8'b00000000 ;
			15'h00000286 : data <= 8'b00000000 ;
			15'h00000287 : data <= 8'b00000000 ;
			15'h00000288 : data <= 8'b00000000 ;
			15'h00000289 : data <= 8'b00000000 ;
			15'h0000028A : data <= 8'b00000000 ;
			15'h0000028B : data <= 8'b00000000 ;
			15'h0000028C : data <= 8'b00000000 ;
			15'h0000028D : data <= 8'b00000000 ;
			15'h0000028E : data <= 8'b00000000 ;
			15'h0000028F : data <= 8'b00000000 ;
			15'h00000290 : data <= 8'b00000000 ;
			15'h00000291 : data <= 8'b00000000 ;
			15'h00000292 : data <= 8'b00000000 ;
			15'h00000293 : data <= 8'b00000000 ;
			15'h00000294 : data <= 8'b00000000 ;
			15'h00000295 : data <= 8'b00000000 ;
			15'h00000296 : data <= 8'b00000000 ;
			15'h00000297 : data <= 8'b00000000 ;
			15'h00000298 : data <= 8'b00000000 ;
			15'h00000299 : data <= 8'b00000000 ;
			15'h0000029A : data <= 8'b00000000 ;
			15'h0000029B : data <= 8'b00000000 ;
			15'h0000029C : data <= 8'b00000000 ;
			15'h0000029D : data <= 8'b00000000 ;
			15'h0000029E : data <= 8'b00000000 ;
			15'h0000029F : data <= 8'b00000000 ;
			15'h000002A0 : data <= 8'b00000000 ;
			15'h000002A1 : data <= 8'b00000000 ;
			15'h000002A2 : data <= 8'b00000000 ;
			15'h000002A3 : data <= 8'b00000000 ;
			15'h000002A4 : data <= 8'b00000000 ;
			15'h000002A5 : data <= 8'b00000000 ;
			15'h000002A6 : data <= 8'b00000000 ;
			15'h000002A7 : data <= 8'b00000000 ;
			15'h000002A8 : data <= 8'b00000000 ;
			15'h000002A9 : data <= 8'b00000000 ;
			15'h000002AA : data <= 8'b00000000 ;
			15'h000002AB : data <= 8'b00000000 ;
			15'h000002AC : data <= 8'b00000000 ;
			15'h000002AD : data <= 8'b00000000 ;
			15'h000002AE : data <= 8'b00000000 ;
			15'h000002AF : data <= 8'b00000000 ;
			15'h000002B0 : data <= 8'b00000000 ;
			15'h000002B1 : data <= 8'b00000000 ;
			15'h000002B2 : data <= 8'b00000000 ;
			15'h000002B3 : data <= 8'b00000000 ;
			15'h000002B4 : data <= 8'b00000000 ;
			15'h000002B5 : data <= 8'b00000000 ;
			15'h000002B6 : data <= 8'b00000000 ;
			15'h000002B7 : data <= 8'b00000000 ;
			15'h000002B8 : data <= 8'b00000000 ;
			15'h000002B9 : data <= 8'b00000000 ;
			15'h000002BA : data <= 8'b00000000 ;
			15'h000002BB : data <= 8'b00000000 ;
			15'h000002BC : data <= 8'b00000000 ;
			15'h000002BD : data <= 8'b00000000 ;
			15'h000002BE : data <= 8'b00000000 ;
			15'h000002BF : data <= 8'b00000000 ;
			15'h000002C0 : data <= 8'b00000000 ;
			15'h000002C1 : data <= 8'b00000000 ;
			15'h000002C2 : data <= 8'b00000000 ;
			15'h000002C3 : data <= 8'b00000000 ;
			15'h000002C4 : data <= 8'b00000000 ;
			15'h000002C5 : data <= 8'b00000000 ;
			15'h000002C6 : data <= 8'b00000000 ;
			15'h000002C7 : data <= 8'b00000000 ;
			15'h000002C8 : data <= 8'b00000000 ;
			15'h000002C9 : data <= 8'b00000000 ;
			15'h000002CA : data <= 8'b00000000 ;
			15'h000002CB : data <= 8'b00000000 ;
			15'h000002CC : data <= 8'b00000000 ;
			15'h000002CD : data <= 8'b00000000 ;
			15'h000002CE : data <= 8'b00000000 ;
			15'h000002CF : data <= 8'b00000000 ;
			15'h000002D0 : data <= 8'b00000000 ;
			15'h000002D1 : data <= 8'b00000000 ;
			15'h000002D2 : data <= 8'b00000000 ;
			15'h000002D3 : data <= 8'b00000000 ;
			15'h000002D4 : data <= 8'b00000000 ;
			15'h000002D5 : data <= 8'b00000000 ;
			15'h000002D6 : data <= 8'b00000000 ;
			15'h000002D7 : data <= 8'b00000000 ;
			15'h000002D8 : data <= 8'b00000000 ;
			15'h000002D9 : data <= 8'b00000000 ;
			15'h000002DA : data <= 8'b00000000 ;
			15'h000002DB : data <= 8'b00000000 ;
			15'h000002DC : data <= 8'b00000000 ;
			15'h000002DD : data <= 8'b00000000 ;
			15'h000002DE : data <= 8'b00000000 ;
			15'h000002DF : data <= 8'b00000000 ;
			15'h000002E0 : data <= 8'b00000000 ;
			15'h000002E1 : data <= 8'b00000000 ;
			15'h000002E2 : data <= 8'b00000000 ;
			15'h000002E3 : data <= 8'b00000000 ;
			15'h000002E4 : data <= 8'b00000000 ;
			15'h000002E5 : data <= 8'b00000000 ;
			15'h000002E6 : data <= 8'b00000000 ;
			15'h000002E7 : data <= 8'b00000000 ;
			15'h000002E8 : data <= 8'b00000000 ;
			15'h000002E9 : data <= 8'b00000000 ;
			15'h000002EA : data <= 8'b00000000 ;
			15'h000002EB : data <= 8'b00000000 ;
			15'h000002EC : data <= 8'b00000000 ;
			15'h000002ED : data <= 8'b00000000 ;
			15'h000002EE : data <= 8'b00000000 ;
			15'h000002EF : data <= 8'b00000000 ;
			15'h000002F0 : data <= 8'b00000000 ;
			15'h000002F1 : data <= 8'b00000000 ;
			15'h000002F2 : data <= 8'b00000000 ;
			15'h000002F3 : data <= 8'b00000000 ;
			15'h000002F4 : data <= 8'b00000000 ;
			15'h000002F5 : data <= 8'b00000000 ;
			15'h000002F6 : data <= 8'b00000000 ;
			15'h000002F7 : data <= 8'b00000000 ;
			15'h000002F8 : data <= 8'b00000000 ;
			15'h000002F9 : data <= 8'b00000000 ;
			15'h000002FA : data <= 8'b00000000 ;
			15'h000002FB : data <= 8'b00000000 ;
			15'h000002FC : data <= 8'b00000000 ;
			15'h000002FD : data <= 8'b00000000 ;
			15'h000002FE : data <= 8'b00000000 ;
			15'h000002FF : data <= 8'b00000000 ;
			15'h00000300 : data <= 8'b00000000 ;
			15'h00000301 : data <= 8'b00000000 ;
			15'h00000302 : data <= 8'b00000000 ;
			15'h00000303 : data <= 8'b00000000 ;
			15'h00000304 : data <= 8'b00000000 ;
			15'h00000305 : data <= 8'b00000000 ;
			15'h00000306 : data <= 8'b00000000 ;
			15'h00000307 : data <= 8'b00000000 ;
			15'h00000308 : data <= 8'b00000000 ;
			15'h00000309 : data <= 8'b00000000 ;
			15'h0000030A : data <= 8'b00000000 ;
			15'h0000030B : data <= 8'b00000000 ;
			15'h0000030C : data <= 8'b00000000 ;
			15'h0000030D : data <= 8'b00000000 ;
			15'h0000030E : data <= 8'b00000000 ;
			15'h0000030F : data <= 8'b00000000 ;
			15'h00000310 : data <= 8'b00000000 ;
			15'h00000311 : data <= 8'b00000000 ;
			15'h00000312 : data <= 8'b00000000 ;
			15'h00000313 : data <= 8'b00000000 ;
			15'h00000314 : data <= 8'b00000000 ;
			15'h00000315 : data <= 8'b00000000 ;
			15'h00000316 : data <= 8'b00000000 ;
			15'h00000317 : data <= 8'b00000000 ;
			15'h00000318 : data <= 8'b00000000 ;
			15'h00000319 : data <= 8'b00000000 ;
			15'h0000031A : data <= 8'b00000000 ;
			15'h0000031B : data <= 8'b00000000 ;
			15'h0000031C : data <= 8'b00000000 ;
			15'h0000031D : data <= 8'b00000000 ;
			15'h0000031E : data <= 8'b00000000 ;
			15'h0000031F : data <= 8'b00000000 ;
			15'h00000320 : data <= 8'b00000000 ;
			15'h00000321 : data <= 8'b00000000 ;
			15'h00000322 : data <= 8'b00000000 ;
			15'h00000323 : data <= 8'b00000000 ;
			15'h00000324 : data <= 8'b00000000 ;
			15'h00000325 : data <= 8'b00000000 ;
			15'h00000326 : data <= 8'b00000000 ;
			15'h00000327 : data <= 8'b00000000 ;
			15'h00000328 : data <= 8'b00000000 ;
			15'h00000329 : data <= 8'b00000000 ;
			15'h0000032A : data <= 8'b00000000 ;
			15'h0000032B : data <= 8'b00000000 ;
			15'h0000032C : data <= 8'b00000000 ;
			15'h0000032D : data <= 8'b00000000 ;
			15'h0000032E : data <= 8'b00000000 ;
			15'h0000032F : data <= 8'b00000000 ;
			15'h00000330 : data <= 8'b00000000 ;
			15'h00000331 : data <= 8'b00000000 ;
			15'h00000332 : data <= 8'b00000000 ;
			15'h00000333 : data <= 8'b00000000 ;
			15'h00000334 : data <= 8'b00000000 ;
			15'h00000335 : data <= 8'b00000000 ;
			15'h00000336 : data <= 8'b00000000 ;
			15'h00000337 : data <= 8'b00000000 ;
			15'h00000338 : data <= 8'b00000000 ;
			15'h00000339 : data <= 8'b00000000 ;
			15'h0000033A : data <= 8'b00000000 ;
			15'h0000033B : data <= 8'b00000000 ;
			15'h0000033C : data <= 8'b00000000 ;
			15'h0000033D : data <= 8'b00000000 ;
			15'h0000033E : data <= 8'b00000000 ;
			15'h0000033F : data <= 8'b00000000 ;
			15'h00000340 : data <= 8'b00000000 ;
			15'h00000341 : data <= 8'b00000000 ;
			15'h00000342 : data <= 8'b00000000 ;
			15'h00000343 : data <= 8'b00000000 ;
			15'h00000344 : data <= 8'b00000000 ;
			15'h00000345 : data <= 8'b00000000 ;
			15'h00000346 : data <= 8'b00000000 ;
			15'h00000347 : data <= 8'b00000000 ;
			15'h00000348 : data <= 8'b00000000 ;
			15'h00000349 : data <= 8'b00000000 ;
			15'h0000034A : data <= 8'b00000000 ;
			15'h0000034B : data <= 8'b00000000 ;
			15'h0000034C : data <= 8'b00000000 ;
			15'h0000034D : data <= 8'b00000000 ;
			15'h0000034E : data <= 8'b00000000 ;
			15'h0000034F : data <= 8'b00000000 ;
			15'h00000350 : data <= 8'b00000000 ;
			15'h00000351 : data <= 8'b00000000 ;
			15'h00000352 : data <= 8'b00000000 ;
			15'h00000353 : data <= 8'b00000000 ;
			15'h00000354 : data <= 8'b00000000 ;
			15'h00000355 : data <= 8'b00000000 ;
			15'h00000356 : data <= 8'b00000000 ;
			15'h00000357 : data <= 8'b00000000 ;
			15'h00000358 : data <= 8'b00000000 ;
			15'h00000359 : data <= 8'b00000000 ;
			15'h0000035A : data <= 8'b00000000 ;
			15'h0000035B : data <= 8'b00000000 ;
			15'h0000035C : data <= 8'b00000000 ;
			15'h0000035D : data <= 8'b00000000 ;
			15'h0000035E : data <= 8'b00000000 ;
			15'h0000035F : data <= 8'b00000000 ;
			15'h00000360 : data <= 8'b00000000 ;
			15'h00000361 : data <= 8'b00000000 ;
			15'h00000362 : data <= 8'b00000000 ;
			15'h00000363 : data <= 8'b00000000 ;
			15'h00000364 : data <= 8'b00000000 ;
			15'h00000365 : data <= 8'b00000000 ;
			15'h00000366 : data <= 8'b00000000 ;
			15'h00000367 : data <= 8'b00000000 ;
			15'h00000368 : data <= 8'b00000000 ;
			15'h00000369 : data <= 8'b00000000 ;
			15'h0000036A : data <= 8'b00000000 ;
			15'h0000036B : data <= 8'b00000000 ;
			15'h0000036C : data <= 8'b00000000 ;
			15'h0000036D : data <= 8'b00000000 ;
			15'h0000036E : data <= 8'b00000000 ;
			15'h0000036F : data <= 8'b00000000 ;
			15'h00000370 : data <= 8'b00000000 ;
			15'h00000371 : data <= 8'b00000000 ;
			15'h00000372 : data <= 8'b00000000 ;
			15'h00000373 : data <= 8'b00000000 ;
			15'h00000374 : data <= 8'b00000000 ;
			15'h00000375 : data <= 8'b00000000 ;
			15'h00000376 : data <= 8'b00000000 ;
			15'h00000377 : data <= 8'b00000000 ;
			15'h00000378 : data <= 8'b00000000 ;
			15'h00000379 : data <= 8'b00000000 ;
			15'h0000037A : data <= 8'b00000000 ;
			15'h0000037B : data <= 8'b00000000 ;
			15'h0000037C : data <= 8'b00000000 ;
			15'h0000037D : data <= 8'b00000000 ;
			15'h0000037E : data <= 8'b00000000 ;
			15'h0000037F : data <= 8'b00000000 ;
			15'h00000380 : data <= 8'b00000000 ;
			15'h00000381 : data <= 8'b00000000 ;
			15'h00000382 : data <= 8'b00000000 ;
			15'h00000383 : data <= 8'b00000000 ;
			15'h00000384 : data <= 8'b00000000 ;
			15'h00000385 : data <= 8'b00000000 ;
			15'h00000386 : data <= 8'b00000000 ;
			15'h00000387 : data <= 8'b00000000 ;
			15'h00000388 : data <= 8'b00000000 ;
			15'h00000389 : data <= 8'b00000000 ;
			15'h0000038A : data <= 8'b00000000 ;
			15'h0000038B : data <= 8'b00000000 ;
			15'h0000038C : data <= 8'b00000000 ;
			15'h0000038D : data <= 8'b00000000 ;
			15'h0000038E : data <= 8'b00000000 ;
			15'h0000038F : data <= 8'b00000000 ;
			15'h00000390 : data <= 8'b00000000 ;
			15'h00000391 : data <= 8'b00000000 ;
			15'h00000392 : data <= 8'b00000000 ;
			15'h00000393 : data <= 8'b00000000 ;
			15'h00000394 : data <= 8'b00000000 ;
			15'h00000395 : data <= 8'b00000000 ;
			15'h00000396 : data <= 8'b00000000 ;
			15'h00000397 : data <= 8'b00000000 ;
			15'h00000398 : data <= 8'b00000000 ;
			15'h00000399 : data <= 8'b00000000 ;
			15'h0000039A : data <= 8'b00000000 ;
			15'h0000039B : data <= 8'b00000000 ;
			15'h0000039C : data <= 8'b00000000 ;
			15'h0000039D : data <= 8'b00000000 ;
			15'h0000039E : data <= 8'b00000000 ;
			15'h0000039F : data <= 8'b00000000 ;
			15'h000003A0 : data <= 8'b00000000 ;
			15'h000003A1 : data <= 8'b00000000 ;
			15'h000003A2 : data <= 8'b00000000 ;
			15'h000003A3 : data <= 8'b00000000 ;
			15'h000003A4 : data <= 8'b00000000 ;
			15'h000003A5 : data <= 8'b00000000 ;
			15'h000003A6 : data <= 8'b00000000 ;
			15'h000003A7 : data <= 8'b00000000 ;
			15'h000003A8 : data <= 8'b00000000 ;
			15'h000003A9 : data <= 8'b00000000 ;
			15'h000003AA : data <= 8'b00000000 ;
			15'h000003AB : data <= 8'b00000000 ;
			15'h000003AC : data <= 8'b00000000 ;
			15'h000003AD : data <= 8'b00000000 ;
			15'h000003AE : data <= 8'b00000000 ;
			15'h000003AF : data <= 8'b00000000 ;
			15'h000003B0 : data <= 8'b00000000 ;
			15'h000003B1 : data <= 8'b00000000 ;
			15'h000003B2 : data <= 8'b00000000 ;
			15'h000003B3 : data <= 8'b00000000 ;
			15'h000003B4 : data <= 8'b00000000 ;
			15'h000003B5 : data <= 8'b00000000 ;
			15'h000003B6 : data <= 8'b00000000 ;
			15'h000003B7 : data <= 8'b00000000 ;
			15'h000003B8 : data <= 8'b00000000 ;
			15'h000003B9 : data <= 8'b00000000 ;
			15'h000003BA : data <= 8'b00000000 ;
			15'h000003BB : data <= 8'b00000000 ;
			15'h000003BC : data <= 8'b00000000 ;
			15'h000003BD : data <= 8'b00000000 ;
			15'h000003BE : data <= 8'b00000000 ;
			15'h000003BF : data <= 8'b00000000 ;
			15'h000003C0 : data <= 8'b00000000 ;
			15'h000003C1 : data <= 8'b00000000 ;
			15'h000003C2 : data <= 8'b00000000 ;
			15'h000003C3 : data <= 8'b00000000 ;
			15'h000003C4 : data <= 8'b00000000 ;
			15'h000003C5 : data <= 8'b00000000 ;
			15'h000003C6 : data <= 8'b00000000 ;
			15'h000003C7 : data <= 8'b00000000 ;
			15'h000003C8 : data <= 8'b00000000 ;
			15'h000003C9 : data <= 8'b00000000 ;
			15'h000003CA : data <= 8'b00000000 ;
			15'h000003CB : data <= 8'b00000000 ;
			15'h000003CC : data <= 8'b00000000 ;
			15'h000003CD : data <= 8'b00000000 ;
			15'h000003CE : data <= 8'b00000000 ;
			15'h000003CF : data <= 8'b00000000 ;
			15'h000003D0 : data <= 8'b00000000 ;
			15'h000003D1 : data <= 8'b00000000 ;
			15'h000003D2 : data <= 8'b00000000 ;
			15'h000003D3 : data <= 8'b00000000 ;
			15'h000003D4 : data <= 8'b00000000 ;
			15'h000003D5 : data <= 8'b00000000 ;
			15'h000003D6 : data <= 8'b00000000 ;
			15'h000003D7 : data <= 8'b00000000 ;
			15'h000003D8 : data <= 8'b00000000 ;
			15'h000003D9 : data <= 8'b00000000 ;
			15'h000003DA : data <= 8'b00000000 ;
			15'h000003DB : data <= 8'b00000000 ;
			15'h000003DC : data <= 8'b00000000 ;
			15'h000003DD : data <= 8'b00000000 ;
			15'h000003DE : data <= 8'b00000000 ;
			15'h000003DF : data <= 8'b00000000 ;
			15'h000003E0 : data <= 8'b00000000 ;
			15'h000003E1 : data <= 8'b00000000 ;
			15'h000003E2 : data <= 8'b00000000 ;
			15'h000003E3 : data <= 8'b00000000 ;
			15'h000003E4 : data <= 8'b00000000 ;
			15'h000003E5 : data <= 8'b00000000 ;
			15'h000003E6 : data <= 8'b00000000 ;
			15'h000003E7 : data <= 8'b00000000 ;
			15'h000003E8 : data <= 8'b00000000 ;
			15'h000003E9 : data <= 8'b00000000 ;
			15'h000003EA : data <= 8'b00000000 ;
			15'h000003EB : data <= 8'b00000000 ;
			15'h000003EC : data <= 8'b00000000 ;
			15'h000003ED : data <= 8'b00000000 ;
			15'h000003EE : data <= 8'b00000000 ;
			15'h000003EF : data <= 8'b00000000 ;
			15'h000003F0 : data <= 8'b00000000 ;
			15'h000003F1 : data <= 8'b00000000 ;
			15'h000003F2 : data <= 8'b00000000 ;
			15'h000003F3 : data <= 8'b00000000 ;
			15'h000003F4 : data <= 8'b00000000 ;
			15'h000003F5 : data <= 8'b00000000 ;
			15'h000003F6 : data <= 8'b00000000 ;
			15'h000003F7 : data <= 8'b00000000 ;
			15'h000003F8 : data <= 8'b00000000 ;
			15'h000003F9 : data <= 8'b00000000 ;
			15'h000003FA : data <= 8'b00000000 ;
			15'h000003FB : data <= 8'b00000000 ;
			15'h000003FC : data <= 8'b00000000 ;
			15'h000003FD : data <= 8'b00000000 ;
			15'h000003FE : data <= 8'b00000000 ;
			15'h000003FF : data <= 8'b00000000 ;
			15'h00000400 : data <= 8'b00000000 ;
			15'h00000401 : data <= 8'b00000000 ;
			15'h00000402 : data <= 8'b00000000 ;
			15'h00000403 : data <= 8'b00000000 ;
			15'h00000404 : data <= 8'b00000000 ;
			15'h00000405 : data <= 8'b00000000 ;
			15'h00000406 : data <= 8'b00000000 ;
			15'h00000407 : data <= 8'b00000000 ;
			15'h00000408 : data <= 8'b00000000 ;
			15'h00000409 : data <= 8'b00000000 ;
			15'h0000040A : data <= 8'b00000000 ;
			15'h0000040B : data <= 8'b00000000 ;
			15'h0000040C : data <= 8'b00000000 ;
			15'h0000040D : data <= 8'b00000000 ;
			15'h0000040E : data <= 8'b00000000 ;
			15'h0000040F : data <= 8'b00000000 ;
			15'h00000410 : data <= 8'b00000000 ;
			15'h00000411 : data <= 8'b00000000 ;
			15'h00000412 : data <= 8'b00000000 ;
			15'h00000413 : data <= 8'b00000000 ;
			15'h00000414 : data <= 8'b00000000 ;
			15'h00000415 : data <= 8'b00000000 ;
			15'h00000416 : data <= 8'b00000000 ;
			15'h00000417 : data <= 8'b00000000 ;
			15'h00000418 : data <= 8'b00000000 ;
			15'h00000419 : data <= 8'b00000000 ;
			15'h0000041A : data <= 8'b00000000 ;
			15'h0000041B : data <= 8'b00000000 ;
			15'h0000041C : data <= 8'b00000000 ;
			15'h0000041D : data <= 8'b00000000 ;
			15'h0000041E : data <= 8'b00000000 ;
			15'h0000041F : data <= 8'b00000000 ;
			15'h00000420 : data <= 8'b00000000 ;
			15'h00000421 : data <= 8'b00000000 ;
			15'h00000422 : data <= 8'b00000000 ;
			15'h00000423 : data <= 8'b00000000 ;
			15'h00000424 : data <= 8'b00000000 ;
			15'h00000425 : data <= 8'b00000000 ;
			15'h00000426 : data <= 8'b00000000 ;
			15'h00000427 : data <= 8'b00000000 ;
			15'h00000428 : data <= 8'b00000000 ;
			15'h00000429 : data <= 8'b00000000 ;
			15'h0000042A : data <= 8'b00000000 ;
			15'h0000042B : data <= 8'b00000000 ;
			15'h0000042C : data <= 8'b00000000 ;
			15'h0000042D : data <= 8'b00000000 ;
			15'h0000042E : data <= 8'b00000000 ;
			15'h0000042F : data <= 8'b00000000 ;
			15'h00000430 : data <= 8'b00000000 ;
			15'h00000431 : data <= 8'b00000000 ;
			15'h00000432 : data <= 8'b00000000 ;
			15'h00000433 : data <= 8'b00000000 ;
			15'h00000434 : data <= 8'b00000000 ;
			15'h00000435 : data <= 8'b00000000 ;
			15'h00000436 : data <= 8'b00000000 ;
			15'h00000437 : data <= 8'b00000000 ;
			15'h00000438 : data <= 8'b00000000 ;
			15'h00000439 : data <= 8'b00000000 ;
			15'h0000043A : data <= 8'b00000000 ;
			15'h0000043B : data <= 8'b00000000 ;
			15'h0000043C : data <= 8'b00000000 ;
			15'h0000043D : data <= 8'b00000000 ;
			15'h0000043E : data <= 8'b00000000 ;
			15'h0000043F : data <= 8'b00000000 ;
			15'h00000440 : data <= 8'b00000000 ;
			15'h00000441 : data <= 8'b00000000 ;
			15'h00000442 : data <= 8'b00000000 ;
			15'h00000443 : data <= 8'b00000000 ;
			15'h00000444 : data <= 8'b00000000 ;
			15'h00000445 : data <= 8'b00000000 ;
			15'h00000446 : data <= 8'b00000000 ;
			15'h00000447 : data <= 8'b00000000 ;
			15'h00000448 : data <= 8'b00000000 ;
			15'h00000449 : data <= 8'b00000000 ;
			15'h0000044A : data <= 8'b00000000 ;
			15'h0000044B : data <= 8'b00000000 ;
			15'h0000044C : data <= 8'b00000000 ;
			15'h0000044D : data <= 8'b00000000 ;
			15'h0000044E : data <= 8'b00000000 ;
			15'h0000044F : data <= 8'b00000000 ;
			15'h00000450 : data <= 8'b00000000 ;
			15'h00000451 : data <= 8'b00000000 ;
			15'h00000452 : data <= 8'b00000000 ;
			15'h00000453 : data <= 8'b00000000 ;
			15'h00000454 : data <= 8'b00000000 ;
			15'h00000455 : data <= 8'b00000000 ;
			15'h00000456 : data <= 8'b00000000 ;
			15'h00000457 : data <= 8'b00000000 ;
			15'h00000458 : data <= 8'b00000000 ;
			15'h00000459 : data <= 8'b00000000 ;
			15'h0000045A : data <= 8'b00000000 ;
			15'h0000045B : data <= 8'b00000000 ;
			15'h0000045C : data <= 8'b00000000 ;
			15'h0000045D : data <= 8'b00000000 ;
			15'h0000045E : data <= 8'b00000000 ;
			15'h0000045F : data <= 8'b00000000 ;
			15'h00000460 : data <= 8'b00000000 ;
			15'h00000461 : data <= 8'b00000000 ;
			15'h00000462 : data <= 8'b00000000 ;
			15'h00000463 : data <= 8'b00000000 ;
			15'h00000464 : data <= 8'b00000000 ;
			15'h00000465 : data <= 8'b00000000 ;
			15'h00000466 : data <= 8'b00000000 ;
			15'h00000467 : data <= 8'b00000000 ;
			15'h00000468 : data <= 8'b00000000 ;
			15'h00000469 : data <= 8'b00000000 ;
			15'h0000046A : data <= 8'b00000000 ;
			15'h0000046B : data <= 8'b00000000 ;
			15'h0000046C : data <= 8'b00000000 ;
			15'h0000046D : data <= 8'b00000000 ;
			15'h0000046E : data <= 8'b00000000 ;
			15'h0000046F : data <= 8'b00000000 ;
			15'h00000470 : data <= 8'b00000000 ;
			15'h00000471 : data <= 8'b00000000 ;
			15'h00000472 : data <= 8'b00000000 ;
			15'h00000473 : data <= 8'b00000000 ;
			15'h00000474 : data <= 8'b00000000 ;
			15'h00000475 : data <= 8'b00000000 ;
			15'h00000476 : data <= 8'b00000000 ;
			15'h00000477 : data <= 8'b00000000 ;
			15'h00000478 : data <= 8'b00000000 ;
			15'h00000479 : data <= 8'b00000000 ;
			15'h0000047A : data <= 8'b00000000 ;
			15'h0000047B : data <= 8'b00000000 ;
			15'h0000047C : data <= 8'b00000000 ;
			15'h0000047D : data <= 8'b00000000 ;
			15'h0000047E : data <= 8'b00000000 ;
			15'h0000047F : data <= 8'b00000000 ;
			15'h00000480 : data <= 8'b00000000 ;
			15'h00000481 : data <= 8'b00000000 ;
			15'h00000482 : data <= 8'b00000000 ;
			15'h00000483 : data <= 8'b00000000 ;
			15'h00000484 : data <= 8'b00000000 ;
			15'h00000485 : data <= 8'b00000000 ;
			15'h00000486 : data <= 8'b00000000 ;
			15'h00000487 : data <= 8'b00000000 ;
			15'h00000488 : data <= 8'b00000000 ;
			15'h00000489 : data <= 8'b00000000 ;
			15'h0000048A : data <= 8'b00000000 ;
			15'h0000048B : data <= 8'b00000000 ;
			15'h0000048C : data <= 8'b00000000 ;
			15'h0000048D : data <= 8'b00000000 ;
			15'h0000048E : data <= 8'b00000000 ;
			15'h0000048F : data <= 8'b00000000 ;
			15'h00000490 : data <= 8'b00000000 ;
			15'h00000491 : data <= 8'b00000000 ;
			15'h00000492 : data <= 8'b00000000 ;
			15'h00000493 : data <= 8'b00000000 ;
			15'h00000494 : data <= 8'b00000000 ;
			15'h00000495 : data <= 8'b00000000 ;
			15'h00000496 : data <= 8'b00000000 ;
			15'h00000497 : data <= 8'b00000000 ;
			15'h00000498 : data <= 8'b00000000 ;
			15'h00000499 : data <= 8'b00000000 ;
			15'h0000049A : data <= 8'b00000000 ;
			15'h0000049B : data <= 8'b00000000 ;
			15'h0000049C : data <= 8'b00000000 ;
			15'h0000049D : data <= 8'b00000000 ;
			15'h0000049E : data <= 8'b00000000 ;
			15'h0000049F : data <= 8'b00000000 ;
			15'h000004A0 : data <= 8'b00000000 ;
			15'h000004A1 : data <= 8'b00000000 ;
			15'h000004A2 : data <= 8'b00000000 ;
			15'h000004A3 : data <= 8'b00000000 ;
			15'h000004A4 : data <= 8'b00000000 ;
			15'h000004A5 : data <= 8'b00000000 ;
			15'h000004A6 : data <= 8'b00000000 ;
			15'h000004A7 : data <= 8'b00000000 ;
			15'h000004A8 : data <= 8'b00000000 ;
			15'h000004A9 : data <= 8'b00000000 ;
			15'h000004AA : data <= 8'b00000000 ;
			15'h000004AB : data <= 8'b00000000 ;
			15'h000004AC : data <= 8'b00000000 ;
			15'h000004AD : data <= 8'b00000000 ;
			15'h000004AE : data <= 8'b00000000 ;
			15'h000004AF : data <= 8'b00000000 ;
			15'h000004B0 : data <= 8'b00000000 ;
			15'h000004B1 : data <= 8'b00000000 ;
			15'h000004B2 : data <= 8'b00000000 ;
			15'h000004B3 : data <= 8'b00000000 ;
			15'h000004B4 : data <= 8'b00000000 ;
			15'h000004B5 : data <= 8'b00000000 ;
			15'h000004B6 : data <= 8'b00000000 ;
			15'h000004B7 : data <= 8'b00000000 ;
			15'h000004B8 : data <= 8'b00000000 ;
			15'h000004B9 : data <= 8'b00000000 ;
			15'h000004BA : data <= 8'b00000000 ;
			15'h000004BB : data <= 8'b00000000 ;
			15'h000004BC : data <= 8'b00000000 ;
			15'h000004BD : data <= 8'b00000000 ;
			15'h000004BE : data <= 8'b00000000 ;
			15'h000004BF : data <= 8'b00000000 ;
			15'h000004C0 : data <= 8'b00000000 ;
			15'h000004C1 : data <= 8'b00000000 ;
			15'h000004C2 : data <= 8'b00000000 ;
			15'h000004C3 : data <= 8'b00000000 ;
			15'h000004C4 : data <= 8'b00000000 ;
			15'h000004C5 : data <= 8'b00000000 ;
			15'h000004C6 : data <= 8'b00000000 ;
			15'h000004C7 : data <= 8'b00000000 ;
			15'h000004C8 : data <= 8'b00000000 ;
			15'h000004C9 : data <= 8'b00000000 ;
			15'h000004CA : data <= 8'b00000000 ;
			15'h000004CB : data <= 8'b00000000 ;
			15'h000004CC : data <= 8'b00000000 ;
			15'h000004CD : data <= 8'b00000000 ;
			15'h000004CE : data <= 8'b00000000 ;
			15'h000004CF : data <= 8'b00000000 ;
			15'h000004D0 : data <= 8'b00000000 ;
			15'h000004D1 : data <= 8'b00000000 ;
			15'h000004D2 : data <= 8'b00000000 ;
			15'h000004D3 : data <= 8'b00000000 ;
			15'h000004D4 : data <= 8'b00000000 ;
			15'h000004D5 : data <= 8'b00000000 ;
			15'h000004D6 : data <= 8'b00000000 ;
			15'h000004D7 : data <= 8'b00000000 ;
			15'h000004D8 : data <= 8'b00000000 ;
			15'h000004D9 : data <= 8'b00000000 ;
			15'h000004DA : data <= 8'b00000000 ;
			15'h000004DB : data <= 8'b00000000 ;
			15'h000004DC : data <= 8'b00000000 ;
			15'h000004DD : data <= 8'b00000000 ;
			15'h000004DE : data <= 8'b00000000 ;
			15'h000004DF : data <= 8'b00000000 ;
			15'h000004E0 : data <= 8'b00000000 ;
			15'h000004E1 : data <= 8'b00000000 ;
			15'h000004E2 : data <= 8'b00000000 ;
			15'h000004E3 : data <= 8'b00000000 ;
			15'h000004E4 : data <= 8'b00000000 ;
			15'h000004E5 : data <= 8'b00000000 ;
			15'h000004E6 : data <= 8'b00000000 ;
			15'h000004E7 : data <= 8'b00000000 ;
			15'h000004E8 : data <= 8'b00000000 ;
			15'h000004E9 : data <= 8'b00000000 ;
			15'h000004EA : data <= 8'b00000000 ;
			15'h000004EB : data <= 8'b00000000 ;
			15'h000004EC : data <= 8'b00000000 ;
			15'h000004ED : data <= 8'b00000000 ;
			15'h000004EE : data <= 8'b00000000 ;
			15'h000004EF : data <= 8'b00000000 ;
			15'h000004F0 : data <= 8'b00000000 ;
			15'h000004F1 : data <= 8'b00000000 ;
			15'h000004F2 : data <= 8'b00000000 ;
			15'h000004F3 : data <= 8'b00000000 ;
			15'h000004F4 : data <= 8'b00000000 ;
			15'h000004F5 : data <= 8'b00000000 ;
			15'h000004F6 : data <= 8'b00000000 ;
			15'h000004F7 : data <= 8'b00000000 ;
			15'h000004F8 : data <= 8'b00000000 ;
			15'h000004F9 : data <= 8'b00000000 ;
			15'h000004FA : data <= 8'b00000000 ;
			15'h000004FB : data <= 8'b00000000 ;
			15'h000004FC : data <= 8'b00000000 ;
			15'h000004FD : data <= 8'b00000000 ;
			15'h000004FE : data <= 8'b00000000 ;
			15'h000004FF : data <= 8'b00000000 ;
			15'h00000500 : data <= 8'b00000000 ;
			15'h00000501 : data <= 8'b00000000 ;
			15'h00000502 : data <= 8'b00000000 ;
			15'h00000503 : data <= 8'b00000000 ;
			15'h00000504 : data <= 8'b00000000 ;
			15'h00000505 : data <= 8'b00000000 ;
			15'h00000506 : data <= 8'b00000000 ;
			15'h00000507 : data <= 8'b00000000 ;
			15'h00000508 : data <= 8'b00000000 ;
			15'h00000509 : data <= 8'b00000000 ;
			15'h0000050A : data <= 8'b00000000 ;
			15'h0000050B : data <= 8'b00000000 ;
			15'h0000050C : data <= 8'b00000000 ;
			15'h0000050D : data <= 8'b00000000 ;
			15'h0000050E : data <= 8'b00000000 ;
			15'h0000050F : data <= 8'b00000000 ;
			15'h00000510 : data <= 8'b00000000 ;
			15'h00000511 : data <= 8'b00000000 ;
			15'h00000512 : data <= 8'b00000000 ;
			15'h00000513 : data <= 8'b00000000 ;
			15'h00000514 : data <= 8'b00000000 ;
			15'h00000515 : data <= 8'b00000000 ;
			15'h00000516 : data <= 8'b00000000 ;
			15'h00000517 : data <= 8'b00000000 ;
			15'h00000518 : data <= 8'b00000000 ;
			15'h00000519 : data <= 8'b00000000 ;
			15'h0000051A : data <= 8'b00000000 ;
			15'h0000051B : data <= 8'b00000000 ;
			15'h0000051C : data <= 8'b00000000 ;
			15'h0000051D : data <= 8'b00000000 ;
			15'h0000051E : data <= 8'b00000000 ;
			15'h0000051F : data <= 8'b00000000 ;
			15'h00000520 : data <= 8'b00000000 ;
			15'h00000521 : data <= 8'b00000000 ;
			15'h00000522 : data <= 8'b00000000 ;
			15'h00000523 : data <= 8'b00000000 ;
			15'h00000524 : data <= 8'b00000000 ;
			15'h00000525 : data <= 8'b00000000 ;
			15'h00000526 : data <= 8'b00000000 ;
			15'h00000527 : data <= 8'b00000000 ;
			15'h00000528 : data <= 8'b00000000 ;
			15'h00000529 : data <= 8'b00000000 ;
			15'h0000052A : data <= 8'b00000000 ;
			15'h0000052B : data <= 8'b00000000 ;
			15'h0000052C : data <= 8'b00000000 ;
			15'h0000052D : data <= 8'b00000000 ;
			15'h0000052E : data <= 8'b00000000 ;
			15'h0000052F : data <= 8'b00000000 ;
			15'h00000530 : data <= 8'b00000000 ;
			15'h00000531 : data <= 8'b00000000 ;
			15'h00000532 : data <= 8'b00000000 ;
			15'h00000533 : data <= 8'b00000000 ;
			15'h00000534 : data <= 8'b00000000 ;
			15'h00000535 : data <= 8'b00000000 ;
			15'h00000536 : data <= 8'b00000000 ;
			15'h00000537 : data <= 8'b00000000 ;
			15'h00000538 : data <= 8'b00000000 ;
			15'h00000539 : data <= 8'b00000000 ;
			15'h0000053A : data <= 8'b00000000 ;
			15'h0000053B : data <= 8'b00000000 ;
			15'h0000053C : data <= 8'b00000000 ;
			15'h0000053D : data <= 8'b00000000 ;
			15'h0000053E : data <= 8'b00000000 ;
			15'h0000053F : data <= 8'b00000000 ;
			15'h00000540 : data <= 8'b00000000 ;
			15'h00000541 : data <= 8'b00000000 ;
			15'h00000542 : data <= 8'b00000000 ;
			15'h00000543 : data <= 8'b00000000 ;
			15'h00000544 : data <= 8'b00000000 ;
			15'h00000545 : data <= 8'b00000000 ;
			15'h00000546 : data <= 8'b00000000 ;
			15'h00000547 : data <= 8'b00000000 ;
			15'h00000548 : data <= 8'b00000000 ;
			15'h00000549 : data <= 8'b00000000 ;
			15'h0000054A : data <= 8'b00000000 ;
			15'h0000054B : data <= 8'b00000000 ;
			15'h0000054C : data <= 8'b00000000 ;
			15'h0000054D : data <= 8'b00000000 ;
			15'h0000054E : data <= 8'b00000000 ;
			15'h0000054F : data <= 8'b00000000 ;
			15'h00000550 : data <= 8'b00000000 ;
			15'h00000551 : data <= 8'b00000000 ;
			15'h00000552 : data <= 8'b00000000 ;
			15'h00000553 : data <= 8'b00000000 ;
			15'h00000554 : data <= 8'b00000000 ;
			15'h00000555 : data <= 8'b00000000 ;
			15'h00000556 : data <= 8'b00000000 ;
			15'h00000557 : data <= 8'b00000000 ;
			15'h00000558 : data <= 8'b00000000 ;
			15'h00000559 : data <= 8'b00000000 ;
			15'h0000055A : data <= 8'b00000000 ;
			15'h0000055B : data <= 8'b00000000 ;
			15'h0000055C : data <= 8'b00000000 ;
			15'h0000055D : data <= 8'b00000000 ;
			15'h0000055E : data <= 8'b00000000 ;
			15'h0000055F : data <= 8'b00000000 ;
			15'h00000560 : data <= 8'b00000000 ;
			15'h00000561 : data <= 8'b00000000 ;
			15'h00000562 : data <= 8'b00000000 ;
			15'h00000563 : data <= 8'b00000000 ;
			15'h00000564 : data <= 8'b00000000 ;
			15'h00000565 : data <= 8'b00000000 ;
			15'h00000566 : data <= 8'b00000000 ;
			15'h00000567 : data <= 8'b00000000 ;
			15'h00000568 : data <= 8'b00000000 ;
			15'h00000569 : data <= 8'b00000000 ;
			15'h0000056A : data <= 8'b00000000 ;
			15'h0000056B : data <= 8'b00000000 ;
			15'h0000056C : data <= 8'b00000000 ;
			15'h0000056D : data <= 8'b00000000 ;
			15'h0000056E : data <= 8'b00000000 ;
			15'h0000056F : data <= 8'b00000000 ;
			15'h00000570 : data <= 8'b00000000 ;
			15'h00000571 : data <= 8'b00000000 ;
			15'h00000572 : data <= 8'b00000000 ;
			15'h00000573 : data <= 8'b00000000 ;
			15'h00000574 : data <= 8'b00000000 ;
			15'h00000575 : data <= 8'b00000000 ;
			15'h00000576 : data <= 8'b00000000 ;
			15'h00000577 : data <= 8'b00000000 ;
			15'h00000578 : data <= 8'b00000000 ;
			15'h00000579 : data <= 8'b00000000 ;
			15'h0000057A : data <= 8'b00000000 ;
			15'h0000057B : data <= 8'b00000000 ;
			15'h0000057C : data <= 8'b00000000 ;
			15'h0000057D : data <= 8'b00000000 ;
			15'h0000057E : data <= 8'b00000000 ;
			15'h0000057F : data <= 8'b00000000 ;
			15'h00000580 : data <= 8'b00000000 ;
			15'h00000581 : data <= 8'b00000000 ;
			15'h00000582 : data <= 8'b00000000 ;
			15'h00000583 : data <= 8'b00000000 ;
			15'h00000584 : data <= 8'b00000000 ;
			15'h00000585 : data <= 8'b00000000 ;
			15'h00000586 : data <= 8'b00000000 ;
			15'h00000587 : data <= 8'b00000000 ;
			15'h00000588 : data <= 8'b00000000 ;
			15'h00000589 : data <= 8'b00000000 ;
			15'h0000058A : data <= 8'b00000000 ;
			15'h0000058B : data <= 8'b00000000 ;
			15'h0000058C : data <= 8'b00000000 ;
			15'h0000058D : data <= 8'b00000000 ;
			15'h0000058E : data <= 8'b00000000 ;
			15'h0000058F : data <= 8'b00000000 ;
			15'h00000590 : data <= 8'b00000000 ;
			15'h00000591 : data <= 8'b00000000 ;
			15'h00000592 : data <= 8'b00000000 ;
			15'h00000593 : data <= 8'b00000000 ;
			15'h00000594 : data <= 8'b00000000 ;
			15'h00000595 : data <= 8'b00000000 ;
			15'h00000596 : data <= 8'b00000000 ;
			15'h00000597 : data <= 8'b00000000 ;
			15'h00000598 : data <= 8'b00000000 ;
			15'h00000599 : data <= 8'b00000000 ;
			15'h0000059A : data <= 8'b00000000 ;
			15'h0000059B : data <= 8'b00000000 ;
			15'h0000059C : data <= 8'b00000000 ;
			15'h0000059D : data <= 8'b00000000 ;
			15'h0000059E : data <= 8'b00000000 ;
			15'h0000059F : data <= 8'b00000000 ;
			15'h000005A0 : data <= 8'b00000000 ;
			15'h000005A1 : data <= 8'b00000000 ;
			15'h000005A2 : data <= 8'b00000000 ;
			15'h000005A3 : data <= 8'b00000000 ;
			15'h000005A4 : data <= 8'b00000000 ;
			15'h000005A5 : data <= 8'b00000000 ;
			15'h000005A6 : data <= 8'b00000000 ;
			15'h000005A7 : data <= 8'b00000000 ;
			15'h000005A8 : data <= 8'b00000000 ;
			15'h000005A9 : data <= 8'b00000000 ;
			15'h000005AA : data <= 8'b00000000 ;
			15'h000005AB : data <= 8'b00000000 ;
			15'h000005AC : data <= 8'b00000000 ;
			15'h000005AD : data <= 8'b00000000 ;
			15'h000005AE : data <= 8'b00000000 ;
			15'h000005AF : data <= 8'b00000000 ;
			15'h000005B0 : data <= 8'b00000000 ;
			15'h000005B1 : data <= 8'b00000000 ;
			15'h000005B2 : data <= 8'b00000000 ;
			15'h000005B3 : data <= 8'b00000000 ;
			15'h000005B4 : data <= 8'b00000000 ;
			15'h000005B5 : data <= 8'b00000000 ;
			15'h000005B6 : data <= 8'b00000000 ;
			15'h000005B7 : data <= 8'b00000000 ;
			15'h000005B8 : data <= 8'b00000000 ;
			15'h000005B9 : data <= 8'b00000000 ;
			15'h000005BA : data <= 8'b00000000 ;
			15'h000005BB : data <= 8'b00000000 ;
			15'h000005BC : data <= 8'b00000000 ;
			15'h000005BD : data <= 8'b00000000 ;
			15'h000005BE : data <= 8'b00000000 ;
			15'h000005BF : data <= 8'b00000000 ;
			15'h000005C0 : data <= 8'b00000000 ;
			15'h000005C1 : data <= 8'b00000000 ;
			15'h000005C2 : data <= 8'b00000000 ;
			15'h000005C3 : data <= 8'b00000000 ;
			15'h000005C4 : data <= 8'b00000000 ;
			15'h000005C5 : data <= 8'b00000000 ;
			15'h000005C6 : data <= 8'b00000000 ;
			15'h000005C7 : data <= 8'b00000000 ;
			15'h000005C8 : data <= 8'b00000000 ;
			15'h000005C9 : data <= 8'b00000000 ;
			15'h000005CA : data <= 8'b00000000 ;
			15'h000005CB : data <= 8'b00000000 ;
			15'h000005CC : data <= 8'b00000000 ;
			15'h000005CD : data <= 8'b00000000 ;
			15'h000005CE : data <= 8'b00000000 ;
			15'h000005CF : data <= 8'b00000000 ;
			15'h000005D0 : data <= 8'b00000000 ;
			15'h000005D1 : data <= 8'b00000000 ;
			15'h000005D2 : data <= 8'b00000000 ;
			15'h000005D3 : data <= 8'b00000000 ;
			15'h000005D4 : data <= 8'b00000000 ;
			15'h000005D5 : data <= 8'b00000000 ;
			15'h000005D6 : data <= 8'b00000000 ;
			15'h000005D7 : data <= 8'b00000000 ;
			15'h000005D8 : data <= 8'b00000000 ;
			15'h000005D9 : data <= 8'b00000000 ;
			15'h000005DA : data <= 8'b00000000 ;
			15'h000005DB : data <= 8'b00000000 ;
			15'h000005DC : data <= 8'b00000000 ;
			15'h000005DD : data <= 8'b00000000 ;
			15'h000005DE : data <= 8'b00000000 ;
			15'h000005DF : data <= 8'b00000000 ;
			15'h000005E0 : data <= 8'b00000000 ;
			15'h000005E1 : data <= 8'b00000000 ;
			15'h000005E2 : data <= 8'b00000000 ;
			15'h000005E3 : data <= 8'b00000000 ;
			15'h000005E4 : data <= 8'b00000000 ;
			15'h000005E5 : data <= 8'b00000000 ;
			15'h000005E6 : data <= 8'b00000000 ;
			15'h000005E7 : data <= 8'b00000000 ;
			15'h000005E8 : data <= 8'b00000000 ;
			15'h000005E9 : data <= 8'b00000000 ;
			15'h000005EA : data <= 8'b00000000 ;
			15'h000005EB : data <= 8'b00000000 ;
			15'h000005EC : data <= 8'b00000000 ;
			15'h000005ED : data <= 8'b00000000 ;
			15'h000005EE : data <= 8'b00000000 ;
			15'h000005EF : data <= 8'b00000000 ;
			15'h000005F0 : data <= 8'b00000000 ;
			15'h000005F1 : data <= 8'b00000000 ;
			15'h000005F2 : data <= 8'b00000000 ;
			15'h000005F3 : data <= 8'b00000000 ;
			15'h000005F4 : data <= 8'b00000000 ;
			15'h000005F5 : data <= 8'b00000000 ;
			15'h000005F6 : data <= 8'b00000000 ;
			15'h000005F7 : data <= 8'b00000000 ;
			15'h000005F8 : data <= 8'b00000000 ;
			15'h000005F9 : data <= 8'b00000000 ;
			15'h000005FA : data <= 8'b00000000 ;
			15'h000005FB : data <= 8'b00000000 ;
			15'h000005FC : data <= 8'b00000000 ;
			15'h000005FD : data <= 8'b00000000 ;
			15'h000005FE : data <= 8'b00000000 ;
			15'h000005FF : data <= 8'b00000000 ;
			15'h00000600 : data <= 8'b00000000 ;
			15'h00000601 : data <= 8'b00000000 ;
			15'h00000602 : data <= 8'b00000000 ;
			15'h00000603 : data <= 8'b00000000 ;
			15'h00000604 : data <= 8'b00000000 ;
			15'h00000605 : data <= 8'b00000000 ;
			15'h00000606 : data <= 8'b00000000 ;
			15'h00000607 : data <= 8'b00000000 ;
			15'h00000608 : data <= 8'b00000000 ;
			15'h00000609 : data <= 8'b00000000 ;
			15'h0000060A : data <= 8'b00000000 ;
			15'h0000060B : data <= 8'b00000000 ;
			15'h0000060C : data <= 8'b00000000 ;
			15'h0000060D : data <= 8'b00000000 ;
			15'h0000060E : data <= 8'b00000000 ;
			15'h0000060F : data <= 8'b00000000 ;
			15'h00000610 : data <= 8'b00000000 ;
			15'h00000611 : data <= 8'b00000000 ;
			15'h00000612 : data <= 8'b00000000 ;
			15'h00000613 : data <= 8'b00000000 ;
			15'h00000614 : data <= 8'b00000000 ;
			15'h00000615 : data <= 8'b00000000 ;
			15'h00000616 : data <= 8'b00000000 ;
			15'h00000617 : data <= 8'b00000000 ;
			15'h00000618 : data <= 8'b00000000 ;
			15'h00000619 : data <= 8'b00000000 ;
			15'h0000061A : data <= 8'b00000000 ;
			15'h0000061B : data <= 8'b00000000 ;
			15'h0000061C : data <= 8'b00000000 ;
			15'h0000061D : data <= 8'b00000000 ;
			15'h0000061E : data <= 8'b00000000 ;
			15'h0000061F : data <= 8'b00000000 ;
			15'h00000620 : data <= 8'b00000000 ;
			15'h00000621 : data <= 8'b00000000 ;
			15'h00000622 : data <= 8'b00000000 ;
			15'h00000623 : data <= 8'b00000000 ;
			15'h00000624 : data <= 8'b00000000 ;
			15'h00000625 : data <= 8'b00000000 ;
			15'h00000626 : data <= 8'b00000000 ;
			15'h00000627 : data <= 8'b00000000 ;
			15'h00000628 : data <= 8'b00000000 ;
			15'h00000629 : data <= 8'b00000000 ;
			15'h0000062A : data <= 8'b00000000 ;
			15'h0000062B : data <= 8'b00000000 ;
			15'h0000062C : data <= 8'b00000000 ;
			15'h0000062D : data <= 8'b00000000 ;
			15'h0000062E : data <= 8'b00000000 ;
			15'h0000062F : data <= 8'b00000000 ;
			15'h00000630 : data <= 8'b00000000 ;
			15'h00000631 : data <= 8'b00000000 ;
			15'h00000632 : data <= 8'b00000000 ;
			15'h00000633 : data <= 8'b00000000 ;
			15'h00000634 : data <= 8'b00000000 ;
			15'h00000635 : data <= 8'b00000000 ;
			15'h00000636 : data <= 8'b00000000 ;
			15'h00000637 : data <= 8'b00000000 ;
			15'h00000638 : data <= 8'b00000000 ;
			15'h00000639 : data <= 8'b00000000 ;
			15'h0000063A : data <= 8'b00000000 ;
			15'h0000063B : data <= 8'b00000000 ;
			15'h0000063C : data <= 8'b00000000 ;
			15'h0000063D : data <= 8'b00000000 ;
			15'h0000063E : data <= 8'b00000000 ;
			15'h0000063F : data <= 8'b00000000 ;
			15'h00000640 : data <= 8'b00000000 ;
			15'h00000641 : data <= 8'b00000000 ;
			15'h00000642 : data <= 8'b00000000 ;
			15'h00000643 : data <= 8'b00000000 ;
			15'h00000644 : data <= 8'b00000000 ;
			15'h00000645 : data <= 8'b00000000 ;
			15'h00000646 : data <= 8'b00000000 ;
			15'h00000647 : data <= 8'b00000000 ;
			15'h00000648 : data <= 8'b00000000 ;
			15'h00000649 : data <= 8'b00000000 ;
			15'h0000064A : data <= 8'b00000000 ;
			15'h0000064B : data <= 8'b00000000 ;
			15'h0000064C : data <= 8'b00000000 ;
			15'h0000064D : data <= 8'b00000000 ;
			15'h0000064E : data <= 8'b00000000 ;
			15'h0000064F : data <= 8'b00000000 ;
			15'h00000650 : data <= 8'b00000000 ;
			15'h00000651 : data <= 8'b00000000 ;
			15'h00000652 : data <= 8'b00000000 ;
			15'h00000653 : data <= 8'b00000000 ;
			15'h00000654 : data <= 8'b00000000 ;
			15'h00000655 : data <= 8'b00000000 ;
			15'h00000656 : data <= 8'b00000000 ;
			15'h00000657 : data <= 8'b00000000 ;
			15'h00000658 : data <= 8'b00000000 ;
			15'h00000659 : data <= 8'b00000000 ;
			15'h0000065A : data <= 8'b00000000 ;
			15'h0000065B : data <= 8'b00000000 ;
			15'h0000065C : data <= 8'b00000000 ;
			15'h0000065D : data <= 8'b00000000 ;
			15'h0000065E : data <= 8'b00000000 ;
			15'h0000065F : data <= 8'b00000000 ;
			15'h00000660 : data <= 8'b00000000 ;
			15'h00000661 : data <= 8'b00000000 ;
			15'h00000662 : data <= 8'b00000000 ;
			15'h00000663 : data <= 8'b00000000 ;
			15'h00000664 : data <= 8'b00000000 ;
			15'h00000665 : data <= 8'b00000000 ;
			15'h00000666 : data <= 8'b00000000 ;
			15'h00000667 : data <= 8'b00000000 ;
			15'h00000668 : data <= 8'b00000000 ;
			15'h00000669 : data <= 8'b00000000 ;
			15'h0000066A : data <= 8'b00000000 ;
			15'h0000066B : data <= 8'b00000000 ;
			15'h0000066C : data <= 8'b00000000 ;
			15'h0000066D : data <= 8'b00000000 ;
			15'h0000066E : data <= 8'b00000000 ;
			15'h0000066F : data <= 8'b00000000 ;
			15'h00000670 : data <= 8'b00000000 ;
			15'h00000671 : data <= 8'b00000000 ;
			15'h00000672 : data <= 8'b00000000 ;
			15'h00000673 : data <= 8'b00000000 ;
			15'h00000674 : data <= 8'b00000000 ;
			15'h00000675 : data <= 8'b00000000 ;
			15'h00000676 : data <= 8'b00000000 ;
			15'h00000677 : data <= 8'b00000000 ;
			15'h00000678 : data <= 8'b00000000 ;
			15'h00000679 : data <= 8'b00000000 ;
			15'h0000067A : data <= 8'b00000000 ;
			15'h0000067B : data <= 8'b00000000 ;
			15'h0000067C : data <= 8'b00000000 ;
			15'h0000067D : data <= 8'b00000000 ;
			15'h0000067E : data <= 8'b00000000 ;
			15'h0000067F : data <= 8'b00000000 ;
			15'h00000680 : data <= 8'b00000000 ;
			15'h00000681 : data <= 8'b00000000 ;
			15'h00000682 : data <= 8'b00000000 ;
			15'h00000683 : data <= 8'b00000000 ;
			15'h00000684 : data <= 8'b00000000 ;
			15'h00000685 : data <= 8'b00000000 ;
			15'h00000686 : data <= 8'b00000000 ;
			15'h00000687 : data <= 8'b00000000 ;
			15'h00000688 : data <= 8'b00000000 ;
			15'h00000689 : data <= 8'b00000000 ;
			15'h0000068A : data <= 8'b00000000 ;
			15'h0000068B : data <= 8'b00000000 ;
			15'h0000068C : data <= 8'b00000000 ;
			15'h0000068D : data <= 8'b00000000 ;
			15'h0000068E : data <= 8'b00000000 ;
			15'h0000068F : data <= 8'b00000000 ;
			15'h00000690 : data <= 8'b00000000 ;
			15'h00000691 : data <= 8'b00000000 ;
			15'h00000692 : data <= 8'b00000000 ;
			15'h00000693 : data <= 8'b00000000 ;
			15'h00000694 : data <= 8'b00000000 ;
			15'h00000695 : data <= 8'b00000000 ;
			15'h00000696 : data <= 8'b00000000 ;
			15'h00000697 : data <= 8'b00000000 ;
			15'h00000698 : data <= 8'b00000000 ;
			15'h00000699 : data <= 8'b00000000 ;
			15'h0000069A : data <= 8'b00000000 ;
			15'h0000069B : data <= 8'b00000000 ;
			15'h0000069C : data <= 8'b00000000 ;
			15'h0000069D : data <= 8'b00000000 ;
			15'h0000069E : data <= 8'b00000000 ;
			15'h0000069F : data <= 8'b00000000 ;
			15'h000006A0 : data <= 8'b00000000 ;
			15'h000006A1 : data <= 8'b00000000 ;
			15'h000006A2 : data <= 8'b00000000 ;
			15'h000006A3 : data <= 8'b00000000 ;
			15'h000006A4 : data <= 8'b00000000 ;
			15'h000006A5 : data <= 8'b00000000 ;
			15'h000006A6 : data <= 8'b00000000 ;
			15'h000006A7 : data <= 8'b00000000 ;
			15'h000006A8 : data <= 8'b00000000 ;
			15'h000006A9 : data <= 8'b00000000 ;
			15'h000006AA : data <= 8'b00000000 ;
			15'h000006AB : data <= 8'b00000000 ;
			15'h000006AC : data <= 8'b00000000 ;
			15'h000006AD : data <= 8'b00000000 ;
			15'h000006AE : data <= 8'b00000000 ;
			15'h000006AF : data <= 8'b00000000 ;
			15'h000006B0 : data <= 8'b00000000 ;
			15'h000006B1 : data <= 8'b00000000 ;
			15'h000006B2 : data <= 8'b00000000 ;
			15'h000006B3 : data <= 8'b00000000 ;
			15'h000006B4 : data <= 8'b00000000 ;
			15'h000006B5 : data <= 8'b00000000 ;
			15'h000006B6 : data <= 8'b00000000 ;
			15'h000006B7 : data <= 8'b00000000 ;
			15'h000006B8 : data <= 8'b00000000 ;
			15'h000006B9 : data <= 8'b00000000 ;
			15'h000006BA : data <= 8'b00000000 ;
			15'h000006BB : data <= 8'b00000000 ;
			15'h000006BC : data <= 8'b00000000 ;
			15'h000006BD : data <= 8'b00000000 ;
			15'h000006BE : data <= 8'b00000000 ;
			15'h000006BF : data <= 8'b00000000 ;
			15'h000006C0 : data <= 8'b00000000 ;
			15'h000006C1 : data <= 8'b00000000 ;
			15'h000006C2 : data <= 8'b00000000 ;
			15'h000006C3 : data <= 8'b00000000 ;
			15'h000006C4 : data <= 8'b00000000 ;
			15'h000006C5 : data <= 8'b00000000 ;
			15'h000006C6 : data <= 8'b00000000 ;
			15'h000006C7 : data <= 8'b00000000 ;
			15'h000006C8 : data <= 8'b00000000 ;
			15'h000006C9 : data <= 8'b00000000 ;
			15'h000006CA : data <= 8'b00000000 ;
			15'h000006CB : data <= 8'b00000000 ;
			15'h000006CC : data <= 8'b00000000 ;
			15'h000006CD : data <= 8'b00000000 ;
			15'h000006CE : data <= 8'b00000000 ;
			15'h000006CF : data <= 8'b00000000 ;
			15'h000006D0 : data <= 8'b00000000 ;
			15'h000006D1 : data <= 8'b00000000 ;
			15'h000006D2 : data <= 8'b00000000 ;
			15'h000006D3 : data <= 8'b00000000 ;
			15'h000006D4 : data <= 8'b00000000 ;
			15'h000006D5 : data <= 8'b00000000 ;
			15'h000006D6 : data <= 8'b00000000 ;
			15'h000006D7 : data <= 8'b00000000 ;
			15'h000006D8 : data <= 8'b00000000 ;
			15'h000006D9 : data <= 8'b00000000 ;
			15'h000006DA : data <= 8'b00000000 ;
			15'h000006DB : data <= 8'b00000000 ;
			15'h000006DC : data <= 8'b00000000 ;
			15'h000006DD : data <= 8'b00000000 ;
			15'h000006DE : data <= 8'b00000000 ;
			15'h000006DF : data <= 8'b00000000 ;
			15'h000006E0 : data <= 8'b00000000 ;
			15'h000006E1 : data <= 8'b00000000 ;
			15'h000006E2 : data <= 8'b00000000 ;
			15'h000006E3 : data <= 8'b00000000 ;
			15'h000006E4 : data <= 8'b00000000 ;
			15'h000006E5 : data <= 8'b00000000 ;
			15'h000006E6 : data <= 8'b00000000 ;
			15'h000006E7 : data <= 8'b00000000 ;
			15'h000006E8 : data <= 8'b00000000 ;
			15'h000006E9 : data <= 8'b00000000 ;
			15'h000006EA : data <= 8'b00000000 ;
			15'h000006EB : data <= 8'b00000000 ;
			15'h000006EC : data <= 8'b00000000 ;
			15'h000006ED : data <= 8'b00000000 ;
			15'h000006EE : data <= 8'b00000000 ;
			15'h000006EF : data <= 8'b00000000 ;
			15'h000006F0 : data <= 8'b00000000 ;
			15'h000006F1 : data <= 8'b00000000 ;
			15'h000006F2 : data <= 8'b00000000 ;
			15'h000006F3 : data <= 8'b00000000 ;
			15'h000006F4 : data <= 8'b00000000 ;
			15'h000006F5 : data <= 8'b00000000 ;
			15'h000006F6 : data <= 8'b00000000 ;
			15'h000006F7 : data <= 8'b00000000 ;
			15'h000006F8 : data <= 8'b00000000 ;
			15'h000006F9 : data <= 8'b00000000 ;
			15'h000006FA : data <= 8'b00000000 ;
			15'h000006FB : data <= 8'b00000000 ;
			15'h000006FC : data <= 8'b00000000 ;
			15'h000006FD : data <= 8'b00000000 ;
			15'h000006FE : data <= 8'b00000000 ;
			15'h000006FF : data <= 8'b00000000 ;
			15'h00000700 : data <= 8'b00000000 ;
			15'h00000701 : data <= 8'b00000000 ;
			15'h00000702 : data <= 8'b00000000 ;
			15'h00000703 : data <= 8'b00000000 ;
			15'h00000704 : data <= 8'b00000000 ;
			15'h00000705 : data <= 8'b00000000 ;
			15'h00000706 : data <= 8'b00000000 ;
			15'h00000707 : data <= 8'b00000000 ;
			15'h00000708 : data <= 8'b00000000 ;
			15'h00000709 : data <= 8'b00000000 ;
			15'h0000070A : data <= 8'b00000000 ;
			15'h0000070B : data <= 8'b00000000 ;
			15'h0000070C : data <= 8'b00000000 ;
			15'h0000070D : data <= 8'b00000000 ;
			15'h0000070E : data <= 8'b00000000 ;
			15'h0000070F : data <= 8'b00000000 ;
			15'h00000710 : data <= 8'b00000000 ;
			15'h00000711 : data <= 8'b00000000 ;
			15'h00000712 : data <= 8'b00000000 ;
			15'h00000713 : data <= 8'b00000000 ;
			15'h00000714 : data <= 8'b00000000 ;
			15'h00000715 : data <= 8'b00000000 ;
			15'h00000716 : data <= 8'b00000000 ;
			15'h00000717 : data <= 8'b00000000 ;
			15'h00000718 : data <= 8'b00000000 ;
			15'h00000719 : data <= 8'b00000000 ;
			15'h0000071A : data <= 8'b00000000 ;
			15'h0000071B : data <= 8'b00000000 ;
			15'h0000071C : data <= 8'b00000000 ;
			15'h0000071D : data <= 8'b00000000 ;
			15'h0000071E : data <= 8'b00000000 ;
			15'h0000071F : data <= 8'b00000000 ;
			15'h00000720 : data <= 8'b00000000 ;
			15'h00000721 : data <= 8'b00000000 ;
			15'h00000722 : data <= 8'b00000000 ;
			15'h00000723 : data <= 8'b00000000 ;
			15'h00000724 : data <= 8'b00000000 ;
			15'h00000725 : data <= 8'b00000000 ;
			15'h00000726 : data <= 8'b00000000 ;
			15'h00000727 : data <= 8'b00000000 ;
			15'h00000728 : data <= 8'b00000000 ;
			15'h00000729 : data <= 8'b00000000 ;
			15'h0000072A : data <= 8'b00000000 ;
			15'h0000072B : data <= 8'b00000000 ;
			15'h0000072C : data <= 8'b00000000 ;
			15'h0000072D : data <= 8'b00000000 ;
			15'h0000072E : data <= 8'b00000000 ;
			15'h0000072F : data <= 8'b00000000 ;
			15'h00000730 : data <= 8'b00000000 ;
			15'h00000731 : data <= 8'b00000000 ;
			15'h00000732 : data <= 8'b00000000 ;
			15'h00000733 : data <= 8'b00000000 ;
			15'h00000734 : data <= 8'b00000000 ;
			15'h00000735 : data <= 8'b00000000 ;
			15'h00000736 : data <= 8'b00000000 ;
			15'h00000737 : data <= 8'b00000000 ;
			15'h00000738 : data <= 8'b00000000 ;
			15'h00000739 : data <= 8'b00000000 ;
			15'h0000073A : data <= 8'b00000000 ;
			15'h0000073B : data <= 8'b00000000 ;
			15'h0000073C : data <= 8'b00000000 ;
			15'h0000073D : data <= 8'b00000000 ;
			15'h0000073E : data <= 8'b00000000 ;
			15'h0000073F : data <= 8'b00000000 ;
			15'h00000740 : data <= 8'b00000000 ;
			15'h00000741 : data <= 8'b00000000 ;
			15'h00000742 : data <= 8'b00000000 ;
			15'h00000743 : data <= 8'b00000000 ;
			15'h00000744 : data <= 8'b00000000 ;
			15'h00000745 : data <= 8'b00000000 ;
			15'h00000746 : data <= 8'b00000000 ;
			15'h00000747 : data <= 8'b00000000 ;
			15'h00000748 : data <= 8'b00000000 ;
			15'h00000749 : data <= 8'b00000000 ;
			15'h0000074A : data <= 8'b00000000 ;
			15'h0000074B : data <= 8'b00000000 ;
			15'h0000074C : data <= 8'b00000000 ;
			15'h0000074D : data <= 8'b00000000 ;
			15'h0000074E : data <= 8'b00000000 ;
			15'h0000074F : data <= 8'b00000000 ;
			15'h00000750 : data <= 8'b00000000 ;
			15'h00000751 : data <= 8'b00000000 ;
			15'h00000752 : data <= 8'b00000000 ;
			15'h00000753 : data <= 8'b00000000 ;
			15'h00000754 : data <= 8'b00000000 ;
			15'h00000755 : data <= 8'b00000000 ;
			15'h00000756 : data <= 8'b00000000 ;
			15'h00000757 : data <= 8'b00000000 ;
			15'h00000758 : data <= 8'b00000000 ;
			15'h00000759 : data <= 8'b00000000 ;
			15'h0000075A : data <= 8'b00000000 ;
			15'h0000075B : data <= 8'b00000000 ;
			15'h0000075C : data <= 8'b00000000 ;
			15'h0000075D : data <= 8'b00000000 ;
			15'h0000075E : data <= 8'b00000000 ;
			15'h0000075F : data <= 8'b00000000 ;
			15'h00000760 : data <= 8'b00000000 ;
			15'h00000761 : data <= 8'b00000000 ;
			15'h00000762 : data <= 8'b00000000 ;
			15'h00000763 : data <= 8'b00000000 ;
			15'h00000764 : data <= 8'b00000000 ;
			15'h00000765 : data <= 8'b00000000 ;
			15'h00000766 : data <= 8'b00000000 ;
			15'h00000767 : data <= 8'b00000000 ;
			15'h00000768 : data <= 8'b00000000 ;
			15'h00000769 : data <= 8'b00000000 ;
			15'h0000076A : data <= 8'b00000000 ;
			15'h0000076B : data <= 8'b00000000 ;
			15'h0000076C : data <= 8'b00000000 ;
			15'h0000076D : data <= 8'b00000000 ;
			15'h0000076E : data <= 8'b00000000 ;
			15'h0000076F : data <= 8'b00000000 ;
			15'h00000770 : data <= 8'b00000000 ;
			15'h00000771 : data <= 8'b00000000 ;
			15'h00000772 : data <= 8'b00000000 ;
			15'h00000773 : data <= 8'b00000000 ;
			15'h00000774 : data <= 8'b00000000 ;
			15'h00000775 : data <= 8'b00000000 ;
			15'h00000776 : data <= 8'b00000000 ;
			15'h00000777 : data <= 8'b00000000 ;
			15'h00000778 : data <= 8'b00000000 ;
			15'h00000779 : data <= 8'b00000000 ;
			15'h0000077A : data <= 8'b00000000 ;
			15'h0000077B : data <= 8'b00000000 ;
			15'h0000077C : data <= 8'b00000000 ;
			15'h0000077D : data <= 8'b00000000 ;
			15'h0000077E : data <= 8'b00000000 ;
			15'h0000077F : data <= 8'b00000000 ;
			15'h00000780 : data <= 8'b00000000 ;
			15'h00000781 : data <= 8'b00000000 ;
			15'h00000782 : data <= 8'b00000000 ;
			15'h00000783 : data <= 8'b00000000 ;
			15'h00000784 : data <= 8'b00000000 ;
			15'h00000785 : data <= 8'b00000000 ;
			15'h00000786 : data <= 8'b00000000 ;
			15'h00000787 : data <= 8'b00000000 ;
			15'h00000788 : data <= 8'b00000000 ;
			15'h00000789 : data <= 8'b00000000 ;
			15'h0000078A : data <= 8'b00000000 ;
			15'h0000078B : data <= 8'b00000000 ;
			15'h0000078C : data <= 8'b00000000 ;
			15'h0000078D : data <= 8'b00000000 ;
			15'h0000078E : data <= 8'b00000000 ;
			15'h0000078F : data <= 8'b00000000 ;
			15'h00000790 : data <= 8'b00000000 ;
			15'h00000791 : data <= 8'b00000000 ;
			15'h00000792 : data <= 8'b00000000 ;
			15'h00000793 : data <= 8'b00000000 ;
			15'h00000794 : data <= 8'b00000000 ;
			15'h00000795 : data <= 8'b00000000 ;
			15'h00000796 : data <= 8'b00000000 ;
			15'h00000797 : data <= 8'b00000000 ;
			15'h00000798 : data <= 8'b00000000 ;
			15'h00000799 : data <= 8'b00000000 ;
			15'h0000079A : data <= 8'b00000000 ;
			15'h0000079B : data <= 8'b00000000 ;
			15'h0000079C : data <= 8'b00000000 ;
			15'h0000079D : data <= 8'b00000000 ;
			15'h0000079E : data <= 8'b00000000 ;
			15'h0000079F : data <= 8'b00000000 ;
			15'h000007A0 : data <= 8'b00000000 ;
			15'h000007A1 : data <= 8'b00000000 ;
			15'h000007A2 : data <= 8'b00000000 ;
			15'h000007A3 : data <= 8'b00000000 ;
			15'h000007A4 : data <= 8'b00000000 ;
			15'h000007A5 : data <= 8'b00000000 ;
			15'h000007A6 : data <= 8'b00000000 ;
			15'h000007A7 : data <= 8'b00000000 ;
			15'h000007A8 : data <= 8'b00000000 ;
			15'h000007A9 : data <= 8'b00000000 ;
			15'h000007AA : data <= 8'b00000000 ;
			15'h000007AB : data <= 8'b00000000 ;
			15'h000007AC : data <= 8'b00000000 ;
			15'h000007AD : data <= 8'b00000000 ;
			15'h000007AE : data <= 8'b00000000 ;
			15'h000007AF : data <= 8'b00000000 ;
			15'h000007B0 : data <= 8'b00000000 ;
			15'h000007B1 : data <= 8'b00000000 ;
			15'h000007B2 : data <= 8'b00000000 ;
			15'h000007B3 : data <= 8'b00000000 ;
			15'h000007B4 : data <= 8'b00000000 ;
			15'h000007B5 : data <= 8'b00000000 ;
			15'h000007B6 : data <= 8'b00000000 ;
			15'h000007B7 : data <= 8'b00000000 ;
			15'h000007B8 : data <= 8'b00000000 ;
			15'h000007B9 : data <= 8'b00000000 ;
			15'h000007BA : data <= 8'b00000000 ;
			15'h000007BB : data <= 8'b00000000 ;
			15'h000007BC : data <= 8'b00000000 ;
			15'h000007BD : data <= 8'b00000000 ;
			15'h000007BE : data <= 8'b00000000 ;
			15'h000007BF : data <= 8'b00000000 ;
			15'h000007C0 : data <= 8'b00000000 ;
			15'h000007C1 : data <= 8'b00000000 ;
			15'h000007C2 : data <= 8'b00000000 ;
			15'h000007C3 : data <= 8'b00000000 ;
			15'h000007C4 : data <= 8'b00000000 ;
			15'h000007C5 : data <= 8'b00000000 ;
			15'h000007C6 : data <= 8'b00000000 ;
			15'h000007C7 : data <= 8'b00000000 ;
			15'h000007C8 : data <= 8'b00000000 ;
			15'h000007C9 : data <= 8'b00000000 ;
			15'h000007CA : data <= 8'b00000000 ;
			15'h000007CB : data <= 8'b00000000 ;
			15'h000007CC : data <= 8'b00000000 ;
			15'h000007CD : data <= 8'b00000000 ;
			15'h000007CE : data <= 8'b00000000 ;
			15'h000007CF : data <= 8'b00000000 ;
			15'h000007D0 : data <= 8'b00000000 ;
			15'h000007D1 : data <= 8'b00000000 ;
			15'h000007D2 : data <= 8'b00000000 ;
			15'h000007D3 : data <= 8'b00000000 ;
			15'h000007D4 : data <= 8'b00000000 ;
			15'h000007D5 : data <= 8'b00000000 ;
			15'h000007D6 : data <= 8'b00000000 ;
			15'h000007D7 : data <= 8'b00000000 ;
			15'h000007D8 : data <= 8'b00000000 ;
			15'h000007D9 : data <= 8'b00000000 ;
			15'h000007DA : data <= 8'b00000000 ;
			15'h000007DB : data <= 8'b00000000 ;
			15'h000007DC : data <= 8'b00000000 ;
			15'h000007DD : data <= 8'b00000000 ;
			15'h000007DE : data <= 8'b00000000 ;
			15'h000007DF : data <= 8'b00000000 ;
			15'h000007E0 : data <= 8'b00000000 ;
			15'h000007E1 : data <= 8'b00000000 ;
			15'h000007E2 : data <= 8'b00000000 ;
			15'h000007E3 : data <= 8'b00000000 ;
			15'h000007E4 : data <= 8'b00000000 ;
			15'h000007E5 : data <= 8'b00000000 ;
			15'h000007E6 : data <= 8'b00000000 ;
			15'h000007E7 : data <= 8'b00000000 ;
			15'h000007E8 : data <= 8'b00000000 ;
			15'h000007E9 : data <= 8'b00000000 ;
			15'h000007EA : data <= 8'b00000000 ;
			15'h000007EB : data <= 8'b00000000 ;
			15'h000007EC : data <= 8'b00000000 ;
			15'h000007ED : data <= 8'b00000000 ;
			15'h000007EE : data <= 8'b00000000 ;
			15'h000007EF : data <= 8'b00000000 ;
			15'h000007F0 : data <= 8'b00000000 ;
			15'h000007F1 : data <= 8'b00000000 ;
			15'h000007F2 : data <= 8'b00000000 ;
			15'h000007F3 : data <= 8'b00000000 ;
			15'h000007F4 : data <= 8'b00000000 ;
			15'h000007F5 : data <= 8'b00000000 ;
			15'h000007F6 : data <= 8'b00000000 ;
			15'h000007F7 : data <= 8'b00000000 ;
			15'h000007F8 : data <= 8'b00000000 ;
			15'h000007F9 : data <= 8'b00000000 ;
			15'h000007FA : data <= 8'b00000000 ;
			15'h000007FB : data <= 8'b00000000 ;
			15'h000007FC : data <= 8'b00000000 ;
			15'h000007FD : data <= 8'b00000000 ;
			15'h000007FE : data <= 8'b00000000 ;
			15'h000007FF : data <= 8'b00000000 ;
			15'h00000800 : data <= 8'b00000000 ;
			15'h00000801 : data <= 8'b00000000 ;
			15'h00000802 : data <= 8'b00000000 ;
			15'h00000803 : data <= 8'b00000000 ;
			15'h00000804 : data <= 8'b00000000 ;
			15'h00000805 : data <= 8'b00000000 ;
			15'h00000806 : data <= 8'b00000000 ;
			15'h00000807 : data <= 8'b00000000 ;
			15'h00000808 : data <= 8'b00000000 ;
			15'h00000809 : data <= 8'b00000000 ;
			15'h0000080A : data <= 8'b00000000 ;
			15'h0000080B : data <= 8'b00000000 ;
			15'h0000080C : data <= 8'b00000000 ;
			15'h0000080D : data <= 8'b00000000 ;
			15'h0000080E : data <= 8'b00000000 ;
			15'h0000080F : data <= 8'b00000000 ;
			15'h00000810 : data <= 8'b00000000 ;
			15'h00000811 : data <= 8'b00000000 ;
			15'h00000812 : data <= 8'b00000000 ;
			15'h00000813 : data <= 8'b00000000 ;
			15'h00000814 : data <= 8'b00000000 ;
			15'h00000815 : data <= 8'b00000000 ;
			15'h00000816 : data <= 8'b00000000 ;
			15'h00000817 : data <= 8'b00000000 ;
			15'h00000818 : data <= 8'b00000000 ;
			15'h00000819 : data <= 8'b00000000 ;
			15'h0000081A : data <= 8'b00000000 ;
			15'h0000081B : data <= 8'b00000000 ;
			15'h0000081C : data <= 8'b00000000 ;
			15'h0000081D : data <= 8'b00000000 ;
			15'h0000081E : data <= 8'b00000000 ;
			15'h0000081F : data <= 8'b00000000 ;
			15'h00000820 : data <= 8'b00000000 ;
			15'h00000821 : data <= 8'b00000000 ;
			15'h00000822 : data <= 8'b00000000 ;
			15'h00000823 : data <= 8'b00000000 ;
			15'h00000824 : data <= 8'b00000000 ;
			15'h00000825 : data <= 8'b00000000 ;
			15'h00000826 : data <= 8'b00000000 ;
			15'h00000827 : data <= 8'b00000000 ;
			15'h00000828 : data <= 8'b00000000 ;
			15'h00000829 : data <= 8'b00000000 ;
			15'h0000082A : data <= 8'b00000000 ;
			15'h0000082B : data <= 8'b00000000 ;
			15'h0000082C : data <= 8'b00000000 ;
			15'h0000082D : data <= 8'b00000000 ;
			15'h0000082E : data <= 8'b00000000 ;
			15'h0000082F : data <= 8'b00000000 ;
			15'h00000830 : data <= 8'b00000000 ;
			15'h00000831 : data <= 8'b00000000 ;
			15'h00000832 : data <= 8'b00000000 ;
			15'h00000833 : data <= 8'b00000000 ;
			15'h00000834 : data <= 8'b00000000 ;
			15'h00000835 : data <= 8'b00000000 ;
			15'h00000836 : data <= 8'b00000000 ;
			15'h00000837 : data <= 8'b00000000 ;
			15'h00000838 : data <= 8'b00000000 ;
			15'h00000839 : data <= 8'b00000000 ;
			15'h0000083A : data <= 8'b00000000 ;
			15'h0000083B : data <= 8'b00000000 ;
			15'h0000083C : data <= 8'b00000000 ;
			15'h0000083D : data <= 8'b00000000 ;
			15'h0000083E : data <= 8'b00000000 ;
			15'h0000083F : data <= 8'b00000000 ;
			15'h00000840 : data <= 8'b00000000 ;
			15'h00000841 : data <= 8'b00000000 ;
			15'h00000842 : data <= 8'b00000000 ;
			15'h00000843 : data <= 8'b00000000 ;
			15'h00000844 : data <= 8'b00000000 ;
			15'h00000845 : data <= 8'b00000000 ;
			15'h00000846 : data <= 8'b00000000 ;
			15'h00000847 : data <= 8'b00000000 ;
			15'h00000848 : data <= 8'b00000000 ;
			15'h00000849 : data <= 8'b00000000 ;
			15'h0000084A : data <= 8'b00000000 ;
			15'h0000084B : data <= 8'b00000000 ;
			15'h0000084C : data <= 8'b00000000 ;
			15'h0000084D : data <= 8'b00000000 ;
			15'h0000084E : data <= 8'b00000000 ;
			15'h0000084F : data <= 8'b00000000 ;
			15'h00000850 : data <= 8'b00000000 ;
			15'h00000851 : data <= 8'b00000000 ;
			15'h00000852 : data <= 8'b00000000 ;
			15'h00000853 : data <= 8'b00000000 ;
			15'h00000854 : data <= 8'b00000000 ;
			15'h00000855 : data <= 8'b00000000 ;
			15'h00000856 : data <= 8'b00000000 ;
			15'h00000857 : data <= 8'b00000000 ;
			15'h00000858 : data <= 8'b00000000 ;
			15'h00000859 : data <= 8'b00000000 ;
			15'h0000085A : data <= 8'b00000000 ;
			15'h0000085B : data <= 8'b00000000 ;
			15'h0000085C : data <= 8'b00000000 ;
			15'h0000085D : data <= 8'b00000000 ;
			15'h0000085E : data <= 8'b00000000 ;
			15'h0000085F : data <= 8'b00000000 ;
			15'h00000860 : data <= 8'b00000000 ;
			15'h00000861 : data <= 8'b00000000 ;
			15'h00000862 : data <= 8'b00000000 ;
			15'h00000863 : data <= 8'b00000000 ;
			15'h00000864 : data <= 8'b00000000 ;
			15'h00000865 : data <= 8'b00000000 ;
			15'h00000866 : data <= 8'b00000000 ;
			15'h00000867 : data <= 8'b00000000 ;
			15'h00000868 : data <= 8'b00000000 ;
			15'h00000869 : data <= 8'b00000000 ;
			15'h0000086A : data <= 8'b00000000 ;
			15'h0000086B : data <= 8'b00000000 ;
			15'h0000086C : data <= 8'b00000000 ;
			15'h0000086D : data <= 8'b00000000 ;
			15'h0000086E : data <= 8'b00000000 ;
			15'h0000086F : data <= 8'b00000000 ;
			15'h00000870 : data <= 8'b00000000 ;
			15'h00000871 : data <= 8'b00000000 ;
			15'h00000872 : data <= 8'b00000000 ;
			15'h00000873 : data <= 8'b00000000 ;
			15'h00000874 : data <= 8'b00000000 ;
			15'h00000875 : data <= 8'b00000000 ;
			15'h00000876 : data <= 8'b00000000 ;
			15'h00000877 : data <= 8'b00000000 ;
			15'h00000878 : data <= 8'b00000000 ;
			15'h00000879 : data <= 8'b00000000 ;
			15'h0000087A : data <= 8'b00000000 ;
			15'h0000087B : data <= 8'b00000000 ;
			15'h0000087C : data <= 8'b00000000 ;
			15'h0000087D : data <= 8'b00000000 ;
			15'h0000087E : data <= 8'b00000000 ;
			15'h0000087F : data <= 8'b00000000 ;
			15'h00000880 : data <= 8'b00000000 ;
			15'h00000881 : data <= 8'b00000000 ;
			15'h00000882 : data <= 8'b00000000 ;
			15'h00000883 : data <= 8'b00000000 ;
			15'h00000884 : data <= 8'b00000000 ;
			15'h00000885 : data <= 8'b00000000 ;
			15'h00000886 : data <= 8'b00000000 ;
			15'h00000887 : data <= 8'b00000000 ;
			15'h00000888 : data <= 8'b00000000 ;
			15'h00000889 : data <= 8'b00000000 ;
			15'h0000088A : data <= 8'b00000000 ;
			15'h0000088B : data <= 8'b00000000 ;
			15'h0000088C : data <= 8'b00000000 ;
			15'h0000088D : data <= 8'b00000000 ;
			15'h0000088E : data <= 8'b00000000 ;
			15'h0000088F : data <= 8'b00000000 ;
			15'h00000890 : data <= 8'b00000000 ;
			15'h00000891 : data <= 8'b00000000 ;
			15'h00000892 : data <= 8'b00000000 ;
			15'h00000893 : data <= 8'b00000000 ;
			15'h00000894 : data <= 8'b00000000 ;
			15'h00000895 : data <= 8'b00000000 ;
			15'h00000896 : data <= 8'b00000000 ;
			15'h00000897 : data <= 8'b00000000 ;
			15'h00000898 : data <= 8'b00000000 ;
			15'h00000899 : data <= 8'b00000000 ;
			15'h0000089A : data <= 8'b00000000 ;
			15'h0000089B : data <= 8'b00000000 ;
			15'h0000089C : data <= 8'b00000000 ;
			15'h0000089D : data <= 8'b00000000 ;
			15'h0000089E : data <= 8'b00000000 ;
			15'h0000089F : data <= 8'b00000000 ;
			15'h000008A0 : data <= 8'b00000000 ;
			15'h000008A1 : data <= 8'b00000000 ;
			15'h000008A2 : data <= 8'b00000000 ;
			15'h000008A3 : data <= 8'b00000000 ;
			15'h000008A4 : data <= 8'b00000000 ;
			15'h000008A5 : data <= 8'b00000000 ;
			15'h000008A6 : data <= 8'b00000000 ;
			15'h000008A7 : data <= 8'b00000000 ;
			15'h000008A8 : data <= 8'b00000000 ;
			15'h000008A9 : data <= 8'b00000000 ;
			15'h000008AA : data <= 8'b00000000 ;
			15'h000008AB : data <= 8'b00000000 ;
			15'h000008AC : data <= 8'b00000000 ;
			15'h000008AD : data <= 8'b00000000 ;
			15'h000008AE : data <= 8'b00000000 ;
			15'h000008AF : data <= 8'b00000000 ;
			15'h000008B0 : data <= 8'b00000000 ;
			15'h000008B1 : data <= 8'b00000000 ;
			15'h000008B2 : data <= 8'b00000000 ;
			15'h000008B3 : data <= 8'b00000000 ;
			15'h000008B4 : data <= 8'b00000000 ;
			15'h000008B5 : data <= 8'b00000000 ;
			15'h000008B6 : data <= 8'b00000000 ;
			15'h000008B7 : data <= 8'b00000000 ;
			15'h000008B8 : data <= 8'b00000000 ;
			15'h000008B9 : data <= 8'b00000000 ;
			15'h000008BA : data <= 8'b00000000 ;
			15'h000008BB : data <= 8'b00000000 ;
			15'h000008BC : data <= 8'b00000000 ;
			15'h000008BD : data <= 8'b00000000 ;
			15'h000008BE : data <= 8'b00000000 ;
			15'h000008BF : data <= 8'b00000000 ;
			15'h000008C0 : data <= 8'b00000000 ;
			15'h000008C1 : data <= 8'b00000000 ;
			15'h000008C2 : data <= 8'b00000000 ;
			15'h000008C3 : data <= 8'b00000000 ;
			15'h000008C4 : data <= 8'b00000000 ;
			15'h000008C5 : data <= 8'b00000000 ;
			15'h000008C6 : data <= 8'b00000000 ;
			15'h000008C7 : data <= 8'b00000000 ;
			15'h000008C8 : data <= 8'b00000000 ;
			15'h000008C9 : data <= 8'b00000000 ;
			15'h000008CA : data <= 8'b00000000 ;
			15'h000008CB : data <= 8'b00000000 ;
			15'h000008CC : data <= 8'b00000000 ;
			15'h000008CD : data <= 8'b00000000 ;
			15'h000008CE : data <= 8'b00000000 ;
			15'h000008CF : data <= 8'b00000000 ;
			15'h000008D0 : data <= 8'b00000000 ;
			15'h000008D1 : data <= 8'b00000000 ;
			15'h000008D2 : data <= 8'b00000000 ;
			15'h000008D3 : data <= 8'b00000000 ;
			15'h000008D4 : data <= 8'b00000000 ;
			15'h000008D5 : data <= 8'b00000000 ;
			15'h000008D6 : data <= 8'b00000000 ;
			15'h000008D7 : data <= 8'b00000000 ;
			15'h000008D8 : data <= 8'b00000000 ;
			15'h000008D9 : data <= 8'b00000000 ;
			15'h000008DA : data <= 8'b00000000 ;
			15'h000008DB : data <= 8'b00000000 ;
			15'h000008DC : data <= 8'b00000000 ;
			15'h000008DD : data <= 8'b00000000 ;
			15'h000008DE : data <= 8'b00000000 ;
			15'h000008DF : data <= 8'b00000000 ;
			15'h000008E0 : data <= 8'b00000000 ;
			15'h000008E1 : data <= 8'b00000000 ;
			15'h000008E2 : data <= 8'b00000000 ;
			15'h000008E3 : data <= 8'b00000000 ;
			15'h000008E4 : data <= 8'b00000000 ;
			15'h000008E5 : data <= 8'b00000000 ;
			15'h000008E6 : data <= 8'b00000000 ;
			15'h000008E7 : data <= 8'b00000000 ;
			15'h000008E8 : data <= 8'b00000000 ;
			15'h000008E9 : data <= 8'b00000000 ;
			15'h000008EA : data <= 8'b00000000 ;
			15'h000008EB : data <= 8'b00000000 ;
			15'h000008EC : data <= 8'b00000000 ;
			15'h000008ED : data <= 8'b00000000 ;
			15'h000008EE : data <= 8'b00000000 ;
			15'h000008EF : data <= 8'b00000000 ;
			15'h000008F0 : data <= 8'b00000000 ;
			15'h000008F1 : data <= 8'b00000000 ;
			15'h000008F2 : data <= 8'b00000000 ;
			15'h000008F3 : data <= 8'b00000000 ;
			15'h000008F4 : data <= 8'b00000000 ;
			15'h000008F5 : data <= 8'b00000000 ;
			15'h000008F6 : data <= 8'b00000000 ;
			15'h000008F7 : data <= 8'b00000000 ;
			15'h000008F8 : data <= 8'b00000000 ;
			15'h000008F9 : data <= 8'b00000000 ;
			15'h000008FA : data <= 8'b00000000 ;
			15'h000008FB : data <= 8'b00000000 ;
			15'h000008FC : data <= 8'b00000000 ;
			15'h000008FD : data <= 8'b00000000 ;
			15'h000008FE : data <= 8'b00000000 ;
			15'h000008FF : data <= 8'b00000000 ;
			15'h00000900 : data <= 8'b00000000 ;
			15'h00000901 : data <= 8'b00000000 ;
			15'h00000902 : data <= 8'b00000000 ;
			15'h00000903 : data <= 8'b00000000 ;
			15'h00000904 : data <= 8'b00000000 ;
			15'h00000905 : data <= 8'b00000000 ;
			15'h00000906 : data <= 8'b00000000 ;
			15'h00000907 : data <= 8'b00000000 ;
			15'h00000908 : data <= 8'b00000000 ;
			15'h00000909 : data <= 8'b00000000 ;
			15'h0000090A : data <= 8'b00000000 ;
			15'h0000090B : data <= 8'b00000000 ;
			15'h0000090C : data <= 8'b00000000 ;
			15'h0000090D : data <= 8'b00000000 ;
			15'h0000090E : data <= 8'b00000000 ;
			15'h0000090F : data <= 8'b00000000 ;
			15'h00000910 : data <= 8'b00000000 ;
			15'h00000911 : data <= 8'b00000000 ;
			15'h00000912 : data <= 8'b00000000 ;
			15'h00000913 : data <= 8'b00000000 ;
			15'h00000914 : data <= 8'b00000000 ;
			15'h00000915 : data <= 8'b00000000 ;
			15'h00000916 : data <= 8'b00000000 ;
			15'h00000917 : data <= 8'b00000000 ;
			15'h00000918 : data <= 8'b00000000 ;
			15'h00000919 : data <= 8'b00000000 ;
			15'h0000091A : data <= 8'b00000000 ;
			15'h0000091B : data <= 8'b00000000 ;
			15'h0000091C : data <= 8'b00000000 ;
			15'h0000091D : data <= 8'b00000000 ;
			15'h0000091E : data <= 8'b00000000 ;
			15'h0000091F : data <= 8'b00000000 ;
			15'h00000920 : data <= 8'b00000000 ;
			15'h00000921 : data <= 8'b00000000 ;
			15'h00000922 : data <= 8'b00000000 ;
			15'h00000923 : data <= 8'b00000000 ;
			15'h00000924 : data <= 8'b00000000 ;
			15'h00000925 : data <= 8'b00000000 ;
			15'h00000926 : data <= 8'b00000000 ;
			15'h00000927 : data <= 8'b00000000 ;
			15'h00000928 : data <= 8'b00000000 ;
			15'h00000929 : data <= 8'b00000000 ;
			15'h0000092A : data <= 8'b00000000 ;
			15'h0000092B : data <= 8'b00000000 ;
			15'h0000092C : data <= 8'b00000000 ;
			15'h0000092D : data <= 8'b00000000 ;
			15'h0000092E : data <= 8'b00000000 ;
			15'h0000092F : data <= 8'b00000000 ;
			15'h00000930 : data <= 8'b00000000 ;
			15'h00000931 : data <= 8'b00000000 ;
			15'h00000932 : data <= 8'b00000000 ;
			15'h00000933 : data <= 8'b00000000 ;
			15'h00000934 : data <= 8'b00000000 ;
			15'h00000935 : data <= 8'b00000000 ;
			15'h00000936 : data <= 8'b00000000 ;
			15'h00000937 : data <= 8'b00000000 ;
			15'h00000938 : data <= 8'b00000000 ;
			15'h00000939 : data <= 8'b00000000 ;
			15'h0000093A : data <= 8'b00000000 ;
			15'h0000093B : data <= 8'b00000000 ;
			15'h0000093C : data <= 8'b00000000 ;
			15'h0000093D : data <= 8'b00000000 ;
			15'h0000093E : data <= 8'b00000000 ;
			15'h0000093F : data <= 8'b00000000 ;
			15'h00000940 : data <= 8'b00000000 ;
			15'h00000941 : data <= 8'b00000000 ;
			15'h00000942 : data <= 8'b00000000 ;
			15'h00000943 : data <= 8'b00000000 ;
			15'h00000944 : data <= 8'b00000000 ;
			15'h00000945 : data <= 8'b00000000 ;
			15'h00000946 : data <= 8'b00000000 ;
			15'h00000947 : data <= 8'b00000000 ;
			15'h00000948 : data <= 8'b00000000 ;
			15'h00000949 : data <= 8'b00000000 ;
			15'h0000094A : data <= 8'b00000000 ;
			15'h0000094B : data <= 8'b00000000 ;
			15'h0000094C : data <= 8'b00000000 ;
			15'h0000094D : data <= 8'b00000000 ;
			15'h0000094E : data <= 8'b00000000 ;
			15'h0000094F : data <= 8'b00000000 ;
			15'h00000950 : data <= 8'b00000000 ;
			15'h00000951 : data <= 8'b00000000 ;
			15'h00000952 : data <= 8'b00000000 ;
			15'h00000953 : data <= 8'b00000000 ;
			15'h00000954 : data <= 8'b00000000 ;
			15'h00000955 : data <= 8'b00000000 ;
			15'h00000956 : data <= 8'b00000000 ;
			15'h00000957 : data <= 8'b00000000 ;
			15'h00000958 : data <= 8'b00000000 ;
			15'h00000959 : data <= 8'b00000000 ;
			15'h0000095A : data <= 8'b00000000 ;
			15'h0000095B : data <= 8'b00000000 ;
			15'h0000095C : data <= 8'b00000000 ;
			15'h0000095D : data <= 8'b00000000 ;
			15'h0000095E : data <= 8'b00000000 ;
			15'h0000095F : data <= 8'b00000000 ;
			15'h00000960 : data <= 8'b00000000 ;
			15'h00000961 : data <= 8'b00000000 ;
			15'h00000962 : data <= 8'b00000000 ;
			15'h00000963 : data <= 8'b00000000 ;
			15'h00000964 : data <= 8'b00000000 ;
			15'h00000965 : data <= 8'b00000000 ;
			15'h00000966 : data <= 8'b00000000 ;
			15'h00000967 : data <= 8'b00000000 ;
			15'h00000968 : data <= 8'b00000000 ;
			15'h00000969 : data <= 8'b00000000 ;
			15'h0000096A : data <= 8'b00000000 ;
			15'h0000096B : data <= 8'b00000000 ;
			15'h0000096C : data <= 8'b00000000 ;
			15'h0000096D : data <= 8'b00000000 ;
			15'h0000096E : data <= 8'b00000000 ;
			15'h0000096F : data <= 8'b00000000 ;
			15'h00000970 : data <= 8'b00000000 ;
			15'h00000971 : data <= 8'b00000000 ;
			15'h00000972 : data <= 8'b00000000 ;
			15'h00000973 : data <= 8'b00000000 ;
			15'h00000974 : data <= 8'b00000000 ;
			15'h00000975 : data <= 8'b00000000 ;
			15'h00000976 : data <= 8'b00000000 ;
			15'h00000977 : data <= 8'b00000000 ;
			15'h00000978 : data <= 8'b00000000 ;
			15'h00000979 : data <= 8'b00000000 ;
			15'h0000097A : data <= 8'b00000000 ;
			15'h0000097B : data <= 8'b00000000 ;
			15'h0000097C : data <= 8'b00000000 ;
			15'h0000097D : data <= 8'b00000000 ;
			15'h0000097E : data <= 8'b00000000 ;
			15'h0000097F : data <= 8'b00000000 ;
			15'h00000980 : data <= 8'b00000000 ;
			15'h00000981 : data <= 8'b00000000 ;
			15'h00000982 : data <= 8'b00000000 ;
			15'h00000983 : data <= 8'b00000000 ;
			15'h00000984 : data <= 8'b00000000 ;
			15'h00000985 : data <= 8'b00000000 ;
			15'h00000986 : data <= 8'b00000000 ;
			15'h00000987 : data <= 8'b00000000 ;
			15'h00000988 : data <= 8'b00000000 ;
			15'h00000989 : data <= 8'b00000000 ;
			15'h0000098A : data <= 8'b00000000 ;
			15'h0000098B : data <= 8'b00000000 ;
			15'h0000098C : data <= 8'b00000000 ;
			15'h0000098D : data <= 8'b00000000 ;
			15'h0000098E : data <= 8'b00000000 ;
			15'h0000098F : data <= 8'b00000000 ;
			15'h00000990 : data <= 8'b00000000 ;
			15'h00000991 : data <= 8'b00000000 ;
			15'h00000992 : data <= 8'b00000000 ;
			15'h00000993 : data <= 8'b00000000 ;
			15'h00000994 : data <= 8'b00000000 ;
			15'h00000995 : data <= 8'b00000000 ;
			15'h00000996 : data <= 8'b00000000 ;
			15'h00000997 : data <= 8'b00000000 ;
			15'h00000998 : data <= 8'b00000000 ;
			15'h00000999 : data <= 8'b00000000 ;
			15'h0000099A : data <= 8'b00000000 ;
			15'h0000099B : data <= 8'b00000000 ;
			15'h0000099C : data <= 8'b00000000 ;
			15'h0000099D : data <= 8'b00000000 ;
			15'h0000099E : data <= 8'b00000000 ;
			15'h0000099F : data <= 8'b00000000 ;
			15'h000009A0 : data <= 8'b00000000 ;
			15'h000009A1 : data <= 8'b00000000 ;
			15'h000009A2 : data <= 8'b00000000 ;
			15'h000009A3 : data <= 8'b00000000 ;
			15'h000009A4 : data <= 8'b00000000 ;
			15'h000009A5 : data <= 8'b00000000 ;
			15'h000009A6 : data <= 8'b00000000 ;
			15'h000009A7 : data <= 8'b00000000 ;
			15'h000009A8 : data <= 8'b00000000 ;
			15'h000009A9 : data <= 8'b00000000 ;
			15'h000009AA : data <= 8'b00000000 ;
			15'h000009AB : data <= 8'b00000000 ;
			15'h000009AC : data <= 8'b00000000 ;
			15'h000009AD : data <= 8'b00000000 ;
			15'h000009AE : data <= 8'b00000000 ;
			15'h000009AF : data <= 8'b00000000 ;
			15'h000009B0 : data <= 8'b00000000 ;
			15'h000009B1 : data <= 8'b00000000 ;
			15'h000009B2 : data <= 8'b00000000 ;
			15'h000009B3 : data <= 8'b00000000 ;
			15'h000009B4 : data <= 8'b00000000 ;
			15'h000009B5 : data <= 8'b00000000 ;
			15'h000009B6 : data <= 8'b00000000 ;
			15'h000009B7 : data <= 8'b00000000 ;
			15'h000009B8 : data <= 8'b00000000 ;
			15'h000009B9 : data <= 8'b00000000 ;
			15'h000009BA : data <= 8'b00000000 ;
			15'h000009BB : data <= 8'b00000000 ;
			15'h000009BC : data <= 8'b00000000 ;
			15'h000009BD : data <= 8'b00000000 ;
			15'h000009BE : data <= 8'b00000000 ;
			15'h000009BF : data <= 8'b00000000 ;
			15'h000009C0 : data <= 8'b00000000 ;
			15'h000009C1 : data <= 8'b00000000 ;
			15'h000009C2 : data <= 8'b00000000 ;
			15'h000009C3 : data <= 8'b00000000 ;
			15'h000009C4 : data <= 8'b00000000 ;
			15'h000009C5 : data <= 8'b00000000 ;
			15'h000009C6 : data <= 8'b00000000 ;
			15'h000009C7 : data <= 8'b00000000 ;
			15'h000009C8 : data <= 8'b00000000 ;
			15'h000009C9 : data <= 8'b00000000 ;
			15'h000009CA : data <= 8'b00000000 ;
			15'h000009CB : data <= 8'b00000000 ;
			15'h000009CC : data <= 8'b00000000 ;
			15'h000009CD : data <= 8'b00000000 ;
			15'h000009CE : data <= 8'b00000000 ;
			15'h000009CF : data <= 8'b00000000 ;
			15'h000009D0 : data <= 8'b00000000 ;
			15'h000009D1 : data <= 8'b00000000 ;
			15'h000009D2 : data <= 8'b00000000 ;
			15'h000009D3 : data <= 8'b00000000 ;
			15'h000009D4 : data <= 8'b00000000 ;
			15'h000009D5 : data <= 8'b00000000 ;
			15'h000009D6 : data <= 8'b00000000 ;
			15'h000009D7 : data <= 8'b00000000 ;
			15'h000009D8 : data <= 8'b00000000 ;
			15'h000009D9 : data <= 8'b00000000 ;
			15'h000009DA : data <= 8'b00000000 ;
			15'h000009DB : data <= 8'b00000000 ;
			15'h000009DC : data <= 8'b00000000 ;
			15'h000009DD : data <= 8'b00000000 ;
			15'h000009DE : data <= 8'b00000000 ;
			15'h000009DF : data <= 8'b00000000 ;
			15'h000009E0 : data <= 8'b00000000 ;
			15'h000009E1 : data <= 8'b00000000 ;
			15'h000009E2 : data <= 8'b00000000 ;
			15'h000009E3 : data <= 8'b00000000 ;
			15'h000009E4 : data <= 8'b00000000 ;
			15'h000009E5 : data <= 8'b00000000 ;
			15'h000009E6 : data <= 8'b00000000 ;
			15'h000009E7 : data <= 8'b00000000 ;
			15'h000009E8 : data <= 8'b00000000 ;
			15'h000009E9 : data <= 8'b00000000 ;
			15'h000009EA : data <= 8'b00000000 ;
			15'h000009EB : data <= 8'b00000000 ;
			15'h000009EC : data <= 8'b00000000 ;
			15'h000009ED : data <= 8'b00000000 ;
			15'h000009EE : data <= 8'b00000000 ;
			15'h000009EF : data <= 8'b00000000 ;
			15'h000009F0 : data <= 8'b00000000 ;
			15'h000009F1 : data <= 8'b00000000 ;
			15'h000009F2 : data <= 8'b00000000 ;
			15'h000009F3 : data <= 8'b00000000 ;
			15'h000009F4 : data <= 8'b00000000 ;
			15'h000009F5 : data <= 8'b00000000 ;
			15'h000009F6 : data <= 8'b00000000 ;
			15'h000009F7 : data <= 8'b00000000 ;
			15'h000009F8 : data <= 8'b00000000 ;
			15'h000009F9 : data <= 8'b00000000 ;
			15'h000009FA : data <= 8'b00000000 ;
			15'h000009FB : data <= 8'b00000000 ;
			15'h000009FC : data <= 8'b00000000 ;
			15'h000009FD : data <= 8'b00000000 ;
			15'h000009FE : data <= 8'b00000000 ;
			15'h000009FF : data <= 8'b00000000 ;
			15'h00000A00 : data <= 8'b00000000 ;
			15'h00000A01 : data <= 8'b00000000 ;
			15'h00000A02 : data <= 8'b00000000 ;
			15'h00000A03 : data <= 8'b00000000 ;
			15'h00000A04 : data <= 8'b00000000 ;
			15'h00000A05 : data <= 8'b00000000 ;
			15'h00000A06 : data <= 8'b00000000 ;
			15'h00000A07 : data <= 8'b00000000 ;
			15'h00000A08 : data <= 8'b00000000 ;
			15'h00000A09 : data <= 8'b00000000 ;
			15'h00000A0A : data <= 8'b00000000 ;
			15'h00000A0B : data <= 8'b00000000 ;
			15'h00000A0C : data <= 8'b00000000 ;
			15'h00000A0D : data <= 8'b00000000 ;
			15'h00000A0E : data <= 8'b00000000 ;
			15'h00000A0F : data <= 8'b00000000 ;
			15'h00000A10 : data <= 8'b00000000 ;
			15'h00000A11 : data <= 8'b00000000 ;
			15'h00000A12 : data <= 8'b00000000 ;
			15'h00000A13 : data <= 8'b00000000 ;
			15'h00000A14 : data <= 8'b00000000 ;
			15'h00000A15 : data <= 8'b00000000 ;
			15'h00000A16 : data <= 8'b00000000 ;
			15'h00000A17 : data <= 8'b00000000 ;
			15'h00000A18 : data <= 8'b00000000 ;
			15'h00000A19 : data <= 8'b00000000 ;
			15'h00000A1A : data <= 8'b00000000 ;
			15'h00000A1B : data <= 8'b00000000 ;
			15'h00000A1C : data <= 8'b00000000 ;
			15'h00000A1D : data <= 8'b00000000 ;
			15'h00000A1E : data <= 8'b00000000 ;
			15'h00000A1F : data <= 8'b00000000 ;
			15'h00000A20 : data <= 8'b00000000 ;
			15'h00000A21 : data <= 8'b00000000 ;
			15'h00000A22 : data <= 8'b00000000 ;
			15'h00000A23 : data <= 8'b00000000 ;
			15'h00000A24 : data <= 8'b00000000 ;
			15'h00000A25 : data <= 8'b00000000 ;
			15'h00000A26 : data <= 8'b00000000 ;
			15'h00000A27 : data <= 8'b00000000 ;
			15'h00000A28 : data <= 8'b00000000 ;
			15'h00000A29 : data <= 8'b00000000 ;
			15'h00000A2A : data <= 8'b00000000 ;
			15'h00000A2B : data <= 8'b00000000 ;
			15'h00000A2C : data <= 8'b00000000 ;
			15'h00000A2D : data <= 8'b00000000 ;
			15'h00000A2E : data <= 8'b00000000 ;
			15'h00000A2F : data <= 8'b00000000 ;
			15'h00000A30 : data <= 8'b00000000 ;
			15'h00000A31 : data <= 8'b00000000 ;
			15'h00000A32 : data <= 8'b00000000 ;
			15'h00000A33 : data <= 8'b00000000 ;
			15'h00000A34 : data <= 8'b00000000 ;
			15'h00000A35 : data <= 8'b00000000 ;
			15'h00000A36 : data <= 8'b00000000 ;
			15'h00000A37 : data <= 8'b00000000 ;
			15'h00000A38 : data <= 8'b00000000 ;
			15'h00000A39 : data <= 8'b00000000 ;
			15'h00000A3A : data <= 8'b00000000 ;
			15'h00000A3B : data <= 8'b00000000 ;
			15'h00000A3C : data <= 8'b00000000 ;
			15'h00000A3D : data <= 8'b00000000 ;
			15'h00000A3E : data <= 8'b00000000 ;
			15'h00000A3F : data <= 8'b00000000 ;
			15'h00000A40 : data <= 8'b00000000 ;
			15'h00000A41 : data <= 8'b00000000 ;
			15'h00000A42 : data <= 8'b00000000 ;
			15'h00000A43 : data <= 8'b00000000 ;
			15'h00000A44 : data <= 8'b00000000 ;
			15'h00000A45 : data <= 8'b00000000 ;
			15'h00000A46 : data <= 8'b00000000 ;
			15'h00000A47 : data <= 8'b00000000 ;
			15'h00000A48 : data <= 8'b00000000 ;
			15'h00000A49 : data <= 8'b00000000 ;
			15'h00000A4A : data <= 8'b00000000 ;
			15'h00000A4B : data <= 8'b00000000 ;
			15'h00000A4C : data <= 8'b00000000 ;
			15'h00000A4D : data <= 8'b00000000 ;
			15'h00000A4E : data <= 8'b00000000 ;
			15'h00000A4F : data <= 8'b00000000 ;
			15'h00000A50 : data <= 8'b00000000 ;
			15'h00000A51 : data <= 8'b00000000 ;
			15'h00000A52 : data <= 8'b00000000 ;
			15'h00000A53 : data <= 8'b00000000 ;
			15'h00000A54 : data <= 8'b00000000 ;
			15'h00000A55 : data <= 8'b00000000 ;
			15'h00000A56 : data <= 8'b00000000 ;
			15'h00000A57 : data <= 8'b00000000 ;
			15'h00000A58 : data <= 8'b00000000 ;
			15'h00000A59 : data <= 8'b00000000 ;
			15'h00000A5A : data <= 8'b00000000 ;
			15'h00000A5B : data <= 8'b00000000 ;
			15'h00000A5C : data <= 8'b00000000 ;
			15'h00000A5D : data <= 8'b00000000 ;
			15'h00000A5E : data <= 8'b00000000 ;
			15'h00000A5F : data <= 8'b00000000 ;
			15'h00000A60 : data <= 8'b00000000 ;
			15'h00000A61 : data <= 8'b00000000 ;
			15'h00000A62 : data <= 8'b00000000 ;
			15'h00000A63 : data <= 8'b00000000 ;
			15'h00000A64 : data <= 8'b00000000 ;
			15'h00000A65 : data <= 8'b00000000 ;
			15'h00000A66 : data <= 8'b00000000 ;
			15'h00000A67 : data <= 8'b00000000 ;
			15'h00000A68 : data <= 8'b00000000 ;
			15'h00000A69 : data <= 8'b00000000 ;
			15'h00000A6A : data <= 8'b00000000 ;
			15'h00000A6B : data <= 8'b00000000 ;
			15'h00000A6C : data <= 8'b00000000 ;
			15'h00000A6D : data <= 8'b00000000 ;
			15'h00000A6E : data <= 8'b00000000 ;
			15'h00000A6F : data <= 8'b00000000 ;
			15'h00000A70 : data <= 8'b00000000 ;
			15'h00000A71 : data <= 8'b00000000 ;
			15'h00000A72 : data <= 8'b00000000 ;
			15'h00000A73 : data <= 8'b00000000 ;
			15'h00000A74 : data <= 8'b00000000 ;
			15'h00000A75 : data <= 8'b00000000 ;
			15'h00000A76 : data <= 8'b00000000 ;
			15'h00000A77 : data <= 8'b00000000 ;
			15'h00000A78 : data <= 8'b00000000 ;
			15'h00000A79 : data <= 8'b00000000 ;
			15'h00000A7A : data <= 8'b00000000 ;
			15'h00000A7B : data <= 8'b00000000 ;
			15'h00000A7C : data <= 8'b00000000 ;
			15'h00000A7D : data <= 8'b00000000 ;
			15'h00000A7E : data <= 8'b00000000 ;
			15'h00000A7F : data <= 8'b00000000 ;
			15'h00000A80 : data <= 8'b00000000 ;
			15'h00000A81 : data <= 8'b00000000 ;
			15'h00000A82 : data <= 8'b00000000 ;
			15'h00000A83 : data <= 8'b00000000 ;
			15'h00000A84 : data <= 8'b00000000 ;
			15'h00000A85 : data <= 8'b00000000 ;
			15'h00000A86 : data <= 8'b00000000 ;
			15'h00000A87 : data <= 8'b00000000 ;
			15'h00000A88 : data <= 8'b00000000 ;
			15'h00000A89 : data <= 8'b00000000 ;
			15'h00000A8A : data <= 8'b00000000 ;
			15'h00000A8B : data <= 8'b00000000 ;
			15'h00000A8C : data <= 8'b00000000 ;
			15'h00000A8D : data <= 8'b00000000 ;
			15'h00000A8E : data <= 8'b00000000 ;
			15'h00000A8F : data <= 8'b00000000 ;
			15'h00000A90 : data <= 8'b00000000 ;
			15'h00000A91 : data <= 8'b00000000 ;
			15'h00000A92 : data <= 8'b00000000 ;
			15'h00000A93 : data <= 8'b00000000 ;
			15'h00000A94 : data <= 8'b00000000 ;
			15'h00000A95 : data <= 8'b00000000 ;
			15'h00000A96 : data <= 8'b00000000 ;
			15'h00000A97 : data <= 8'b00000000 ;
			15'h00000A98 : data <= 8'b00000000 ;
			15'h00000A99 : data <= 8'b00000000 ;
			15'h00000A9A : data <= 8'b00000000 ;
			15'h00000A9B : data <= 8'b00000000 ;
			15'h00000A9C : data <= 8'b00000000 ;
			15'h00000A9D : data <= 8'b00000000 ;
			15'h00000A9E : data <= 8'b00000000 ;
			15'h00000A9F : data <= 8'b00000000 ;
			15'h00000AA0 : data <= 8'b00000000 ;
			15'h00000AA1 : data <= 8'b00000000 ;
			15'h00000AA2 : data <= 8'b00000000 ;
			15'h00000AA3 : data <= 8'b00000000 ;
			15'h00000AA4 : data <= 8'b00000000 ;
			15'h00000AA5 : data <= 8'b00000000 ;
			15'h00000AA6 : data <= 8'b00000000 ;
			15'h00000AA7 : data <= 8'b00000000 ;
			15'h00000AA8 : data <= 8'b00000000 ;
			15'h00000AA9 : data <= 8'b00000000 ;
			15'h00000AAA : data <= 8'b00000000 ;
			15'h00000AAB : data <= 8'b00000000 ;
			15'h00000AAC : data <= 8'b00000000 ;
			15'h00000AAD : data <= 8'b00000000 ;
			15'h00000AAE : data <= 8'b00000000 ;
			15'h00000AAF : data <= 8'b00000000 ;
			15'h00000AB0 : data <= 8'b00000000 ;
			15'h00000AB1 : data <= 8'b00000000 ;
			15'h00000AB2 : data <= 8'b00000000 ;
			15'h00000AB3 : data <= 8'b00000000 ;
			15'h00000AB4 : data <= 8'b00000000 ;
			15'h00000AB5 : data <= 8'b00000000 ;
			15'h00000AB6 : data <= 8'b00000000 ;
			15'h00000AB7 : data <= 8'b00000000 ;
			15'h00000AB8 : data <= 8'b00000000 ;
			15'h00000AB9 : data <= 8'b00000000 ;
			15'h00000ABA : data <= 8'b00000000 ;
			15'h00000ABB : data <= 8'b00000000 ;
			15'h00000ABC : data <= 8'b00000000 ;
			15'h00000ABD : data <= 8'b00000000 ;
			15'h00000ABE : data <= 8'b00000000 ;
			15'h00000ABF : data <= 8'b00000000 ;
			15'h00000AC0 : data <= 8'b00000000 ;
			15'h00000AC1 : data <= 8'b00000000 ;
			15'h00000AC2 : data <= 8'b00000000 ;
			15'h00000AC3 : data <= 8'b00000000 ;
			15'h00000AC4 : data <= 8'b00000000 ;
			15'h00000AC5 : data <= 8'b00000000 ;
			15'h00000AC6 : data <= 8'b00000000 ;
			15'h00000AC7 : data <= 8'b00000000 ;
			15'h00000AC8 : data <= 8'b00000000 ;
			15'h00000AC9 : data <= 8'b00000000 ;
			15'h00000ACA : data <= 8'b00000000 ;
			15'h00000ACB : data <= 8'b00000000 ;
			15'h00000ACC : data <= 8'b00000000 ;
			15'h00000ACD : data <= 8'b00000000 ;
			15'h00000ACE : data <= 8'b00000000 ;
			15'h00000ACF : data <= 8'b00000000 ;
			15'h00000AD0 : data <= 8'b00000000 ;
			15'h00000AD1 : data <= 8'b00000000 ;
			15'h00000AD2 : data <= 8'b00000000 ;
			15'h00000AD3 : data <= 8'b00000000 ;
			15'h00000AD4 : data <= 8'b00000000 ;
			15'h00000AD5 : data <= 8'b00000000 ;
			15'h00000AD6 : data <= 8'b00000000 ;
			15'h00000AD7 : data <= 8'b00000000 ;
			15'h00000AD8 : data <= 8'b00000000 ;
			15'h00000AD9 : data <= 8'b00000000 ;
			15'h00000ADA : data <= 8'b00000000 ;
			15'h00000ADB : data <= 8'b00000000 ;
			15'h00000ADC : data <= 8'b00000000 ;
			15'h00000ADD : data <= 8'b00000000 ;
			15'h00000ADE : data <= 8'b00000000 ;
			15'h00000ADF : data <= 8'b00000000 ;
			15'h00000AE0 : data <= 8'b00000000 ;
			15'h00000AE1 : data <= 8'b00000000 ;
			15'h00000AE2 : data <= 8'b00000000 ;
			15'h00000AE3 : data <= 8'b00000000 ;
			15'h00000AE4 : data <= 8'b00000000 ;
			15'h00000AE5 : data <= 8'b00000000 ;
			15'h00000AE6 : data <= 8'b00000000 ;
			15'h00000AE7 : data <= 8'b00000000 ;
			15'h00000AE8 : data <= 8'b00000000 ;
			15'h00000AE9 : data <= 8'b00000000 ;
			15'h00000AEA : data <= 8'b00000000 ;
			15'h00000AEB : data <= 8'b00000000 ;
			15'h00000AEC : data <= 8'b00000000 ;
			15'h00000AED : data <= 8'b00000000 ;
			15'h00000AEE : data <= 8'b00000000 ;
			15'h00000AEF : data <= 8'b00000000 ;
			15'h00000AF0 : data <= 8'b00000000 ;
			15'h00000AF1 : data <= 8'b00000000 ;
			15'h00000AF2 : data <= 8'b00000000 ;
			15'h00000AF3 : data <= 8'b00000000 ;
			15'h00000AF4 : data <= 8'b00000000 ;
			15'h00000AF5 : data <= 8'b00000000 ;
			15'h00000AF6 : data <= 8'b00000000 ;
			15'h00000AF7 : data <= 8'b00000000 ;
			15'h00000AF8 : data <= 8'b00000000 ;
			15'h00000AF9 : data <= 8'b00000000 ;
			15'h00000AFA : data <= 8'b00000000 ;
			15'h00000AFB : data <= 8'b00000000 ;
			15'h00000AFC : data <= 8'b00000000 ;
			15'h00000AFD : data <= 8'b00000000 ;
			15'h00000AFE : data <= 8'b00000000 ;
			15'h00000AFF : data <= 8'b00000000 ;
			15'h00000B00 : data <= 8'b00000000 ;
			15'h00000B01 : data <= 8'b00000000 ;
			15'h00000B02 : data <= 8'b00000000 ;
			15'h00000B03 : data <= 8'b00000000 ;
			15'h00000B04 : data <= 8'b00000000 ;
			15'h00000B05 : data <= 8'b00000000 ;
			15'h00000B06 : data <= 8'b00000000 ;
			15'h00000B07 : data <= 8'b00000000 ;
			15'h00000B08 : data <= 8'b00000000 ;
			15'h00000B09 : data <= 8'b00000000 ;
			15'h00000B0A : data <= 8'b00000000 ;
			15'h00000B0B : data <= 8'b00000000 ;
			15'h00000B0C : data <= 8'b00000000 ;
			15'h00000B0D : data <= 8'b00000000 ;
			15'h00000B0E : data <= 8'b00000000 ;
			15'h00000B0F : data <= 8'b00000000 ;
			15'h00000B10 : data <= 8'b00000000 ;
			15'h00000B11 : data <= 8'b00000000 ;
			15'h00000B12 : data <= 8'b00000000 ;
			15'h00000B13 : data <= 8'b00000000 ;
			15'h00000B14 : data <= 8'b00000000 ;
			15'h00000B15 : data <= 8'b00000000 ;
			15'h00000B16 : data <= 8'b00000000 ;
			15'h00000B17 : data <= 8'b00000000 ;
			15'h00000B18 : data <= 8'b00000000 ;
			15'h00000B19 : data <= 8'b00000000 ;
			15'h00000B1A : data <= 8'b00000000 ;
			15'h00000B1B : data <= 8'b00000000 ;
			15'h00000B1C : data <= 8'b00000000 ;
			15'h00000B1D : data <= 8'b00000000 ;
			15'h00000B1E : data <= 8'b00000000 ;
			15'h00000B1F : data <= 8'b00000000 ;
			15'h00000B20 : data <= 8'b00000000 ;
			15'h00000B21 : data <= 8'b00000000 ;
			15'h00000B22 : data <= 8'b00000000 ;
			15'h00000B23 : data <= 8'b00000000 ;
			15'h00000B24 : data <= 8'b00000000 ;
			15'h00000B25 : data <= 8'b00000000 ;
			15'h00000B26 : data <= 8'b00000000 ;
			15'h00000B27 : data <= 8'b00000000 ;
			15'h00000B28 : data <= 8'b00000000 ;
			15'h00000B29 : data <= 8'b00000000 ;
			15'h00000B2A : data <= 8'b00000000 ;
			15'h00000B2B : data <= 8'b00000000 ;
			15'h00000B2C : data <= 8'b00000000 ;
			15'h00000B2D : data <= 8'b00000000 ;
			15'h00000B2E : data <= 8'b00000000 ;
			15'h00000B2F : data <= 8'b00000000 ;
			15'h00000B30 : data <= 8'b00000000 ;
			15'h00000B31 : data <= 8'b00000000 ;
			15'h00000B32 : data <= 8'b00000000 ;
			15'h00000B33 : data <= 8'b00000000 ;
			15'h00000B34 : data <= 8'b00000000 ;
			15'h00000B35 : data <= 8'b00000000 ;
			15'h00000B36 : data <= 8'b00000000 ;
			15'h00000B37 : data <= 8'b00000000 ;
			15'h00000B38 : data <= 8'b00000000 ;
			15'h00000B39 : data <= 8'b00000000 ;
			15'h00000B3A : data <= 8'b00000000 ;
			15'h00000B3B : data <= 8'b00000000 ;
			15'h00000B3C : data <= 8'b00000000 ;
			15'h00000B3D : data <= 8'b00000000 ;
			15'h00000B3E : data <= 8'b00000000 ;
			15'h00000B3F : data <= 8'b00000000 ;
			15'h00000B40 : data <= 8'b00000000 ;
			15'h00000B41 : data <= 8'b00000000 ;
			15'h00000B42 : data <= 8'b00000000 ;
			15'h00000B43 : data <= 8'b00000000 ;
			15'h00000B44 : data <= 8'b00000000 ;
			15'h00000B45 : data <= 8'b00000000 ;
			15'h00000B46 : data <= 8'b00000000 ;
			15'h00000B47 : data <= 8'b00000000 ;
			15'h00000B48 : data <= 8'b00000000 ;
			15'h00000B49 : data <= 8'b00000000 ;
			15'h00000B4A : data <= 8'b00000000 ;
			15'h00000B4B : data <= 8'b00000000 ;
			15'h00000B4C : data <= 8'b00000000 ;
			15'h00000B4D : data <= 8'b00000000 ;
			15'h00000B4E : data <= 8'b00000000 ;
			15'h00000B4F : data <= 8'b00000000 ;
			15'h00000B50 : data <= 8'b00000000 ;
			15'h00000B51 : data <= 8'b00000000 ;
			15'h00000B52 : data <= 8'b00000000 ;
			15'h00000B53 : data <= 8'b00000000 ;
			15'h00000B54 : data <= 8'b00000000 ;
			15'h00000B55 : data <= 8'b00000000 ;
			15'h00000B56 : data <= 8'b00000000 ;
			15'h00000B57 : data <= 8'b00000000 ;
			15'h00000B58 : data <= 8'b00000000 ;
			15'h00000B59 : data <= 8'b00000000 ;
			15'h00000B5A : data <= 8'b00000000 ;
			15'h00000B5B : data <= 8'b00000000 ;
			15'h00000B5C : data <= 8'b00000000 ;
			15'h00000B5D : data <= 8'b00000000 ;
			15'h00000B5E : data <= 8'b00000000 ;
			15'h00000B5F : data <= 8'b00000000 ;
			15'h00000B60 : data <= 8'b00000000 ;
			15'h00000B61 : data <= 8'b00000000 ;
			15'h00000B62 : data <= 8'b00000000 ;
			15'h00000B63 : data <= 8'b00000000 ;
			15'h00000B64 : data <= 8'b00000000 ;
			15'h00000B65 : data <= 8'b00000000 ;
			15'h00000B66 : data <= 8'b00000000 ;
			15'h00000B67 : data <= 8'b00000000 ;
			15'h00000B68 : data <= 8'b00000000 ;
			15'h00000B69 : data <= 8'b00000000 ;
			15'h00000B6A : data <= 8'b00000000 ;
			15'h00000B6B : data <= 8'b00000000 ;
			15'h00000B6C : data <= 8'b00000000 ;
			15'h00000B6D : data <= 8'b00000000 ;
			15'h00000B6E : data <= 8'b00000000 ;
			15'h00000B6F : data <= 8'b00000000 ;
			15'h00000B70 : data <= 8'b00000000 ;
			15'h00000B71 : data <= 8'b00000000 ;
			15'h00000B72 : data <= 8'b00000000 ;
			15'h00000B73 : data <= 8'b00000000 ;
			15'h00000B74 : data <= 8'b00000000 ;
			15'h00000B75 : data <= 8'b00000000 ;
			15'h00000B76 : data <= 8'b00000000 ;
			15'h00000B77 : data <= 8'b00000000 ;
			15'h00000B78 : data <= 8'b00000000 ;
			15'h00000B79 : data <= 8'b00000000 ;
			15'h00000B7A : data <= 8'b00000000 ;
			15'h00000B7B : data <= 8'b00000000 ;
			15'h00000B7C : data <= 8'b00000000 ;
			15'h00000B7D : data <= 8'b00000000 ;
			15'h00000B7E : data <= 8'b00000000 ;
			15'h00000B7F : data <= 8'b00000000 ;
			15'h00000B80 : data <= 8'b00000000 ;
			15'h00000B81 : data <= 8'b00000000 ;
			15'h00000B82 : data <= 8'b00000000 ;
			15'h00000B83 : data <= 8'b00000000 ;
			15'h00000B84 : data <= 8'b00000000 ;
			15'h00000B85 : data <= 8'b00000000 ;
			15'h00000B86 : data <= 8'b00000000 ;
			15'h00000B87 : data <= 8'b00000000 ;
			15'h00000B88 : data <= 8'b00000000 ;
			15'h00000B89 : data <= 8'b00000000 ;
			15'h00000B8A : data <= 8'b00000000 ;
			15'h00000B8B : data <= 8'b00000000 ;
			15'h00000B8C : data <= 8'b00000000 ;
			15'h00000B8D : data <= 8'b00000000 ;
			15'h00000B8E : data <= 8'b00000000 ;
			15'h00000B8F : data <= 8'b00000000 ;
			15'h00000B90 : data <= 8'b00000000 ;
			15'h00000B91 : data <= 8'b00000000 ;
			15'h00000B92 : data <= 8'b00000000 ;
			15'h00000B93 : data <= 8'b00000000 ;
			15'h00000B94 : data <= 8'b00000000 ;
			15'h00000B95 : data <= 8'b00000000 ;
			15'h00000B96 : data <= 8'b00000000 ;
			15'h00000B97 : data <= 8'b00000000 ;
			15'h00000B98 : data <= 8'b00000000 ;
			15'h00000B99 : data <= 8'b00000000 ;
			15'h00000B9A : data <= 8'b00000000 ;
			15'h00000B9B : data <= 8'b00000000 ;
			15'h00000B9C : data <= 8'b00000000 ;
			15'h00000B9D : data <= 8'b00000000 ;
			15'h00000B9E : data <= 8'b00000000 ;
			15'h00000B9F : data <= 8'b00000000 ;
			15'h00000BA0 : data <= 8'b00000000 ;
			15'h00000BA1 : data <= 8'b00000000 ;
			15'h00000BA2 : data <= 8'b00000000 ;
			15'h00000BA3 : data <= 8'b00000000 ;
			15'h00000BA4 : data <= 8'b00000000 ;
			15'h00000BA5 : data <= 8'b00000000 ;
			15'h00000BA6 : data <= 8'b00000000 ;
			15'h00000BA7 : data <= 8'b00000000 ;
			15'h00000BA8 : data <= 8'b00000000 ;
			15'h00000BA9 : data <= 8'b00000000 ;
			15'h00000BAA : data <= 8'b00000000 ;
			15'h00000BAB : data <= 8'b00000000 ;
			15'h00000BAC : data <= 8'b00000000 ;
			15'h00000BAD : data <= 8'b00000000 ;
			15'h00000BAE : data <= 8'b00000000 ;
			15'h00000BAF : data <= 8'b00000000 ;
			15'h00000BB0 : data <= 8'b00000000 ;
			15'h00000BB1 : data <= 8'b00000000 ;
			15'h00000BB2 : data <= 8'b00000000 ;
			15'h00000BB3 : data <= 8'b00000000 ;
			15'h00000BB4 : data <= 8'b00000000 ;
			15'h00000BB5 : data <= 8'b00000000 ;
			15'h00000BB6 : data <= 8'b00000000 ;
			15'h00000BB7 : data <= 8'b00000000 ;
			15'h00000BB8 : data <= 8'b00000000 ;
			15'h00000BB9 : data <= 8'b00000000 ;
			15'h00000BBA : data <= 8'b00000000 ;
			15'h00000BBB : data <= 8'b00000000 ;
			15'h00000BBC : data <= 8'b00000000 ;
			15'h00000BBD : data <= 8'b00000000 ;
			15'h00000BBE : data <= 8'b00000000 ;
			15'h00000BBF : data <= 8'b00000000 ;
			15'h00000BC0 : data <= 8'b00000000 ;
			15'h00000BC1 : data <= 8'b00000000 ;
			15'h00000BC2 : data <= 8'b00000000 ;
			15'h00000BC3 : data <= 8'b00000000 ;
			15'h00000BC4 : data <= 8'b00000000 ;
			15'h00000BC5 : data <= 8'b00000000 ;
			15'h00000BC6 : data <= 8'b00000000 ;
			15'h00000BC7 : data <= 8'b00000000 ;
			15'h00000BC8 : data <= 8'b00000000 ;
			15'h00000BC9 : data <= 8'b00000000 ;
			15'h00000BCA : data <= 8'b00000000 ;
			15'h00000BCB : data <= 8'b00000000 ;
			15'h00000BCC : data <= 8'b00000000 ;
			15'h00000BCD : data <= 8'b00000000 ;
			15'h00000BCE : data <= 8'b00000000 ;
			15'h00000BCF : data <= 8'b00000000 ;
			15'h00000BD0 : data <= 8'b00000000 ;
			15'h00000BD1 : data <= 8'b00000000 ;
			15'h00000BD2 : data <= 8'b00000000 ;
			15'h00000BD3 : data <= 8'b00000000 ;
			15'h00000BD4 : data <= 8'b00000000 ;
			15'h00000BD5 : data <= 8'b00000000 ;
			15'h00000BD6 : data <= 8'b00000000 ;
			15'h00000BD7 : data <= 8'b00000000 ;
			15'h00000BD8 : data <= 8'b00000000 ;
			15'h00000BD9 : data <= 8'b00000000 ;
			15'h00000BDA : data <= 8'b00000000 ;
			15'h00000BDB : data <= 8'b00000000 ;
			15'h00000BDC : data <= 8'b00000000 ;
			15'h00000BDD : data <= 8'b00000000 ;
			15'h00000BDE : data <= 8'b00000000 ;
			15'h00000BDF : data <= 8'b00000000 ;
			15'h00000BE0 : data <= 8'b00000000 ;
			15'h00000BE1 : data <= 8'b00000000 ;
			15'h00000BE2 : data <= 8'b00000000 ;
			15'h00000BE3 : data <= 8'b00000000 ;
			15'h00000BE4 : data <= 8'b00000000 ;
			15'h00000BE5 : data <= 8'b00000000 ;
			15'h00000BE6 : data <= 8'b00000000 ;
			15'h00000BE7 : data <= 8'b00000000 ;
			15'h00000BE8 : data <= 8'b00000000 ;
			15'h00000BE9 : data <= 8'b00000000 ;
			15'h00000BEA : data <= 8'b00000000 ;
			15'h00000BEB : data <= 8'b00000000 ;
			15'h00000BEC : data <= 8'b00000000 ;
			15'h00000BED : data <= 8'b00000000 ;
			15'h00000BEE : data <= 8'b00000000 ;
			15'h00000BEF : data <= 8'b00000000 ;
			15'h00000BF0 : data <= 8'b00000000 ;
			15'h00000BF1 : data <= 8'b00000000 ;
			15'h00000BF2 : data <= 8'b00000000 ;
			15'h00000BF3 : data <= 8'b00000000 ;
			15'h00000BF4 : data <= 8'b00000000 ;
			15'h00000BF5 : data <= 8'b00000000 ;
			15'h00000BF6 : data <= 8'b00000000 ;
			15'h00000BF7 : data <= 8'b00000000 ;
			15'h00000BF8 : data <= 8'b00000000 ;
			15'h00000BF9 : data <= 8'b00000000 ;
			15'h00000BFA : data <= 8'b00000000 ;
			15'h00000BFB : data <= 8'b00000000 ;
			15'h00000BFC : data <= 8'b00000000 ;
			15'h00000BFD : data <= 8'b00000000 ;
			15'h00000BFE : data <= 8'b00000000 ;
			15'h00000BFF : data <= 8'b00000000 ;
			15'h00000C00 : data <= 8'b00000000 ;
			15'h00000C01 : data <= 8'b00000000 ;
			15'h00000C02 : data <= 8'b00000000 ;
			15'h00000C03 : data <= 8'b00000000 ;
			15'h00000C04 : data <= 8'b00000000 ;
			15'h00000C05 : data <= 8'b00000000 ;
			15'h00000C06 : data <= 8'b00000000 ;
			15'h00000C07 : data <= 8'b00000000 ;
			15'h00000C08 : data <= 8'b00000000 ;
			15'h00000C09 : data <= 8'b00000000 ;
			15'h00000C0A : data <= 8'b00000000 ;
			15'h00000C0B : data <= 8'b00000000 ;
			15'h00000C0C : data <= 8'b00000000 ;
			15'h00000C0D : data <= 8'b00000000 ;
			15'h00000C0E : data <= 8'b00000000 ;
			15'h00000C0F : data <= 8'b00000000 ;
			15'h00000C10 : data <= 8'b00000000 ;
			15'h00000C11 : data <= 8'b00000000 ;
			15'h00000C12 : data <= 8'b00000000 ;
			15'h00000C13 : data <= 8'b00000000 ;
			15'h00000C14 : data <= 8'b00000000 ;
			15'h00000C15 : data <= 8'b00000000 ;
			15'h00000C16 : data <= 8'b00000000 ;
			15'h00000C17 : data <= 8'b00000000 ;
			15'h00000C18 : data <= 8'b00000000 ;
			15'h00000C19 : data <= 8'b00000000 ;
			15'h00000C1A : data <= 8'b00000000 ;
			15'h00000C1B : data <= 8'b00000000 ;
			15'h00000C1C : data <= 8'b00000000 ;
			15'h00000C1D : data <= 8'b00000000 ;
			15'h00000C1E : data <= 8'b00000000 ;
			15'h00000C1F : data <= 8'b00000000 ;
			15'h00000C20 : data <= 8'b00000000 ;
			15'h00000C21 : data <= 8'b00000000 ;
			15'h00000C22 : data <= 8'b00000000 ;
			15'h00000C23 : data <= 8'b00000000 ;
			15'h00000C24 : data <= 8'b00000000 ;
			15'h00000C25 : data <= 8'b00000000 ;
			15'h00000C26 : data <= 8'b00000000 ;
			15'h00000C27 : data <= 8'b00000000 ;
			15'h00000C28 : data <= 8'b00000000 ;
			15'h00000C29 : data <= 8'b00000000 ;
			15'h00000C2A : data <= 8'b00000000 ;
			15'h00000C2B : data <= 8'b00000000 ;
			15'h00000C2C : data <= 8'b00000000 ;
			15'h00000C2D : data <= 8'b00000000 ;
			15'h00000C2E : data <= 8'b00000000 ;
			15'h00000C2F : data <= 8'b00000000 ;
			15'h00000C30 : data <= 8'b00000000 ;
			15'h00000C31 : data <= 8'b00000000 ;
			15'h00000C32 : data <= 8'b00000000 ;
			15'h00000C33 : data <= 8'b00000000 ;
			15'h00000C34 : data <= 8'b00000000 ;
			15'h00000C35 : data <= 8'b00000000 ;
			15'h00000C36 : data <= 8'b00000000 ;
			15'h00000C37 : data <= 8'b00000000 ;
			15'h00000C38 : data <= 8'b00000000 ;
			15'h00000C39 : data <= 8'b00000000 ;
			15'h00000C3A : data <= 8'b00000000 ;
			15'h00000C3B : data <= 8'b00000000 ;
			15'h00000C3C : data <= 8'b00000000 ;
			15'h00000C3D : data <= 8'b00000000 ;
			15'h00000C3E : data <= 8'b00000000 ;
			15'h00000C3F : data <= 8'b00000000 ;
			15'h00000C40 : data <= 8'b00000000 ;
			15'h00000C41 : data <= 8'b00000000 ;
			15'h00000C42 : data <= 8'b00000000 ;
			15'h00000C43 : data <= 8'b00000000 ;
			15'h00000C44 : data <= 8'b00000000 ;
			15'h00000C45 : data <= 8'b00000000 ;
			15'h00000C46 : data <= 8'b00000000 ;
			15'h00000C47 : data <= 8'b00000000 ;
			15'h00000C48 : data <= 8'b00000000 ;
			15'h00000C49 : data <= 8'b00000000 ;
			15'h00000C4A : data <= 8'b00000000 ;
			15'h00000C4B : data <= 8'b00000000 ;
			15'h00000C4C : data <= 8'b00000000 ;
			15'h00000C4D : data <= 8'b00000000 ;
			15'h00000C4E : data <= 8'b00000000 ;
			15'h00000C4F : data <= 8'b00000000 ;
			15'h00000C50 : data <= 8'b00000000 ;
			15'h00000C51 : data <= 8'b00000000 ;
			15'h00000C52 : data <= 8'b00000000 ;
			15'h00000C53 : data <= 8'b00000000 ;
			15'h00000C54 : data <= 8'b00000000 ;
			15'h00000C55 : data <= 8'b00000000 ;
			15'h00000C56 : data <= 8'b00000000 ;
			15'h00000C57 : data <= 8'b00000000 ;
			15'h00000C58 : data <= 8'b00000000 ;
			15'h00000C59 : data <= 8'b00000000 ;
			15'h00000C5A : data <= 8'b00000000 ;
			15'h00000C5B : data <= 8'b00000000 ;
			15'h00000C5C : data <= 8'b00000000 ;
			15'h00000C5D : data <= 8'b00000000 ;
			15'h00000C5E : data <= 8'b00000000 ;
			15'h00000C5F : data <= 8'b00000000 ;
			15'h00000C60 : data <= 8'b00000000 ;
			15'h00000C61 : data <= 8'b00000000 ;
			15'h00000C62 : data <= 8'b00000000 ;
			15'h00000C63 : data <= 8'b00000000 ;
			15'h00000C64 : data <= 8'b00000000 ;
			15'h00000C65 : data <= 8'b00000000 ;
			15'h00000C66 : data <= 8'b00000000 ;
			15'h00000C67 : data <= 8'b00000000 ;
			15'h00000C68 : data <= 8'b00000000 ;
			15'h00000C69 : data <= 8'b00000000 ;
			15'h00000C6A : data <= 8'b00000000 ;
			15'h00000C6B : data <= 8'b00000000 ;
			15'h00000C6C : data <= 8'b00000000 ;
			15'h00000C6D : data <= 8'b00000000 ;
			15'h00000C6E : data <= 8'b00000000 ;
			15'h00000C6F : data <= 8'b00000000 ;
			15'h00000C70 : data <= 8'b00000000 ;
			15'h00000C71 : data <= 8'b00000000 ;
			15'h00000C72 : data <= 8'b00000000 ;
			15'h00000C73 : data <= 8'b00000000 ;
			15'h00000C74 : data <= 8'b00000000 ;
			15'h00000C75 : data <= 8'b00000000 ;
			15'h00000C76 : data <= 8'b00000000 ;
			15'h00000C77 : data <= 8'b00000000 ;
			15'h00000C78 : data <= 8'b00000000 ;
			15'h00000C79 : data <= 8'b00000000 ;
			15'h00000C7A : data <= 8'b00000000 ;
			15'h00000C7B : data <= 8'b00000000 ;
			15'h00000C7C : data <= 8'b00000000 ;
			15'h00000C7D : data <= 8'b00000000 ;
			15'h00000C7E : data <= 8'b00000000 ;
			15'h00000C7F : data <= 8'b00000000 ;
			15'h00000C80 : data <= 8'b00000000 ;
			15'h00000C81 : data <= 8'b00000000 ;
			15'h00000C82 : data <= 8'b00000000 ;
			15'h00000C83 : data <= 8'b00000000 ;
			15'h00000C84 : data <= 8'b00000000 ;
			15'h00000C85 : data <= 8'b00000000 ;
			15'h00000C86 : data <= 8'b00000000 ;
			15'h00000C87 : data <= 8'b00000000 ;
			15'h00000C88 : data <= 8'b00000000 ;
			15'h00000C89 : data <= 8'b00000000 ;
			15'h00000C8A : data <= 8'b00000000 ;
			15'h00000C8B : data <= 8'b00000000 ;
			15'h00000C8C : data <= 8'b00000000 ;
			15'h00000C8D : data <= 8'b00000000 ;
			15'h00000C8E : data <= 8'b00000000 ;
			15'h00000C8F : data <= 8'b00000000 ;
			15'h00000C90 : data <= 8'b00000000 ;
			15'h00000C91 : data <= 8'b00000000 ;
			15'h00000C92 : data <= 8'b00000000 ;
			15'h00000C93 : data <= 8'b00000000 ;
			15'h00000C94 : data <= 8'b00000000 ;
			15'h00000C95 : data <= 8'b00000000 ;
			15'h00000C96 : data <= 8'b00000000 ;
			15'h00000C97 : data <= 8'b00000000 ;
			15'h00000C98 : data <= 8'b00000000 ;
			15'h00000C99 : data <= 8'b00000000 ;
			15'h00000C9A : data <= 8'b00000000 ;
			15'h00000C9B : data <= 8'b00000000 ;
			15'h00000C9C : data <= 8'b00000000 ;
			15'h00000C9D : data <= 8'b00000000 ;
			15'h00000C9E : data <= 8'b00000000 ;
			15'h00000C9F : data <= 8'b00000000 ;
			15'h00000CA0 : data <= 8'b00000000 ;
			15'h00000CA1 : data <= 8'b00000000 ;
			15'h00000CA2 : data <= 8'b00000000 ;
			15'h00000CA3 : data <= 8'b00000000 ;
			15'h00000CA4 : data <= 8'b00000000 ;
			15'h00000CA5 : data <= 8'b00000000 ;
			15'h00000CA6 : data <= 8'b00000000 ;
			15'h00000CA7 : data <= 8'b00000000 ;
			15'h00000CA8 : data <= 8'b00000000 ;
			15'h00000CA9 : data <= 8'b00000000 ;
			15'h00000CAA : data <= 8'b00000000 ;
			15'h00000CAB : data <= 8'b00000000 ;
			15'h00000CAC : data <= 8'b00000000 ;
			15'h00000CAD : data <= 8'b00000000 ;
			15'h00000CAE : data <= 8'b00000000 ;
			15'h00000CAF : data <= 8'b00000000 ;
			15'h00000CB0 : data <= 8'b00000000 ;
			15'h00000CB1 : data <= 8'b00000000 ;
			15'h00000CB2 : data <= 8'b00000000 ;
			15'h00000CB3 : data <= 8'b00000000 ;
			15'h00000CB4 : data <= 8'b00000000 ;
			15'h00000CB5 : data <= 8'b00000000 ;
			15'h00000CB6 : data <= 8'b00000000 ;
			15'h00000CB7 : data <= 8'b00000000 ;
			15'h00000CB8 : data <= 8'b00000000 ;
			15'h00000CB9 : data <= 8'b00000000 ;
			15'h00000CBA : data <= 8'b00000000 ;
			15'h00000CBB : data <= 8'b00000000 ;
			15'h00000CBC : data <= 8'b00000000 ;
			15'h00000CBD : data <= 8'b00000000 ;
			15'h00000CBE : data <= 8'b00000000 ;
			15'h00000CBF : data <= 8'b00000000 ;
			15'h00000CC0 : data <= 8'b00000000 ;
			15'h00000CC1 : data <= 8'b00000000 ;
			15'h00000CC2 : data <= 8'b00000000 ;
			15'h00000CC3 : data <= 8'b00000000 ;
			15'h00000CC4 : data <= 8'b00000000 ;
			15'h00000CC5 : data <= 8'b00000000 ;
			15'h00000CC6 : data <= 8'b00000000 ;
			15'h00000CC7 : data <= 8'b00000000 ;
			15'h00000CC8 : data <= 8'b00000000 ;
			15'h00000CC9 : data <= 8'b00000000 ;
			15'h00000CCA : data <= 8'b00000000 ;
			15'h00000CCB : data <= 8'b00000000 ;
			15'h00000CCC : data <= 8'b00000000 ;
			15'h00000CCD : data <= 8'b00000000 ;
			15'h00000CCE : data <= 8'b00000000 ;
			15'h00000CCF : data <= 8'b00000000 ;
			15'h00000CD0 : data <= 8'b00000000 ;
			15'h00000CD1 : data <= 8'b00000000 ;
			15'h00000CD2 : data <= 8'b00000000 ;
			15'h00000CD3 : data <= 8'b00000000 ;
			15'h00000CD4 : data <= 8'b00000000 ;
			15'h00000CD5 : data <= 8'b00000000 ;
			15'h00000CD6 : data <= 8'b00000000 ;
			15'h00000CD7 : data <= 8'b00000000 ;
			15'h00000CD8 : data <= 8'b00000000 ;
			15'h00000CD9 : data <= 8'b00000000 ;
			15'h00000CDA : data <= 8'b00000000 ;
			15'h00000CDB : data <= 8'b00000000 ;
			15'h00000CDC : data <= 8'b00000000 ;
			15'h00000CDD : data <= 8'b00000000 ;
			15'h00000CDE : data <= 8'b00000000 ;
			15'h00000CDF : data <= 8'b00000000 ;
			15'h00000CE0 : data <= 8'b00000000 ;
			15'h00000CE1 : data <= 8'b00000000 ;
			15'h00000CE2 : data <= 8'b00000000 ;
			15'h00000CE3 : data <= 8'b00000000 ;
			15'h00000CE4 : data <= 8'b00000000 ;
			15'h00000CE5 : data <= 8'b00000000 ;
			15'h00000CE6 : data <= 8'b00000000 ;
			15'h00000CE7 : data <= 8'b00000000 ;
			15'h00000CE8 : data <= 8'b00000000 ;
			15'h00000CE9 : data <= 8'b00000000 ;
			15'h00000CEA : data <= 8'b00000000 ;
			15'h00000CEB : data <= 8'b00000000 ;
			15'h00000CEC : data <= 8'b00000000 ;
			15'h00000CED : data <= 8'b00000000 ;
			15'h00000CEE : data <= 8'b00000000 ;
			15'h00000CEF : data <= 8'b00000000 ;
			15'h00000CF0 : data <= 8'b00000000 ;
			15'h00000CF1 : data <= 8'b00000000 ;
			15'h00000CF2 : data <= 8'b00000000 ;
			15'h00000CF3 : data <= 8'b00000000 ;
			15'h00000CF4 : data <= 8'b00000000 ;
			15'h00000CF5 : data <= 8'b00000000 ;
			15'h00000CF6 : data <= 8'b00000000 ;
			15'h00000CF7 : data <= 8'b00000000 ;
			15'h00000CF8 : data <= 8'b00000000 ;
			15'h00000CF9 : data <= 8'b00000000 ;
			15'h00000CFA : data <= 8'b00000000 ;
			15'h00000CFB : data <= 8'b00000000 ;
			15'h00000CFC : data <= 8'b00000000 ;
			15'h00000CFD : data <= 8'b00000000 ;
			15'h00000CFE : data <= 8'b00000000 ;
			15'h00000CFF : data <= 8'b00000000 ;
			15'h00000D00 : data <= 8'b00000000 ;
			15'h00000D01 : data <= 8'b00000000 ;
			15'h00000D02 : data <= 8'b00000000 ;
			15'h00000D03 : data <= 8'b00000000 ;
			15'h00000D04 : data <= 8'b00000000 ;
			15'h00000D05 : data <= 8'b00000000 ;
			15'h00000D06 : data <= 8'b00000000 ;
			15'h00000D07 : data <= 8'b00000000 ;
			15'h00000D08 : data <= 8'b00000000 ;
			15'h00000D09 : data <= 8'b00000000 ;
			15'h00000D0A : data <= 8'b00000000 ;
			15'h00000D0B : data <= 8'b00000000 ;
			15'h00000D0C : data <= 8'b00000000 ;
			15'h00000D0D : data <= 8'b00000000 ;
			15'h00000D0E : data <= 8'b00000000 ;
			15'h00000D0F : data <= 8'b00000000 ;
			15'h00000D10 : data <= 8'b00000000 ;
			15'h00000D11 : data <= 8'b00000000 ;
			15'h00000D12 : data <= 8'b00000000 ;
			15'h00000D13 : data <= 8'b00000000 ;
			15'h00000D14 : data <= 8'b00000000 ;
			15'h00000D15 : data <= 8'b00000000 ;
			15'h00000D16 : data <= 8'b00000000 ;
			15'h00000D17 : data <= 8'b00000000 ;
			15'h00000D18 : data <= 8'b00000000 ;
			15'h00000D19 : data <= 8'b00000000 ;
			15'h00000D1A : data <= 8'b00000000 ;
			15'h00000D1B : data <= 8'b00000000 ;
			15'h00000D1C : data <= 8'b00000000 ;
			15'h00000D1D : data <= 8'b00000000 ;
			15'h00000D1E : data <= 8'b00000000 ;
			15'h00000D1F : data <= 8'b00000000 ;
			15'h00000D20 : data <= 8'b00000000 ;
			15'h00000D21 : data <= 8'b00000000 ;
			15'h00000D22 : data <= 8'b00000000 ;
			15'h00000D23 : data <= 8'b00000000 ;
			15'h00000D24 : data <= 8'b00000000 ;
			15'h00000D25 : data <= 8'b00000000 ;
			15'h00000D26 : data <= 8'b00000000 ;
			15'h00000D27 : data <= 8'b00000000 ;
			15'h00000D28 : data <= 8'b00000000 ;
			15'h00000D29 : data <= 8'b00000000 ;
			15'h00000D2A : data <= 8'b00000000 ;
			15'h00000D2B : data <= 8'b00000000 ;
			15'h00000D2C : data <= 8'b00000000 ;
			15'h00000D2D : data <= 8'b00000000 ;
			15'h00000D2E : data <= 8'b00000000 ;
			15'h00000D2F : data <= 8'b00000000 ;
			15'h00000D30 : data <= 8'b00000000 ;
			15'h00000D31 : data <= 8'b00000000 ;
			15'h00000D32 : data <= 8'b00000000 ;
			15'h00000D33 : data <= 8'b00000000 ;
			15'h00000D34 : data <= 8'b00000000 ;
			15'h00000D35 : data <= 8'b00000000 ;
			15'h00000D36 : data <= 8'b00000000 ;
			15'h00000D37 : data <= 8'b00000000 ;
			15'h00000D38 : data <= 8'b00000000 ;
			15'h00000D39 : data <= 8'b00000000 ;
			15'h00000D3A : data <= 8'b00000000 ;
			15'h00000D3B : data <= 8'b00000000 ;
			15'h00000D3C : data <= 8'b00000000 ;
			15'h00000D3D : data <= 8'b00000000 ;
			15'h00000D3E : data <= 8'b00000000 ;
			15'h00000D3F : data <= 8'b00000000 ;
			15'h00000D40 : data <= 8'b00000000 ;
			15'h00000D41 : data <= 8'b00000000 ;
			15'h00000D42 : data <= 8'b00000000 ;
			15'h00000D43 : data <= 8'b00000000 ;
			15'h00000D44 : data <= 8'b00000000 ;
			15'h00000D45 : data <= 8'b00000000 ;
			15'h00000D46 : data <= 8'b00000000 ;
			15'h00000D47 : data <= 8'b00000000 ;
			15'h00000D48 : data <= 8'b00000000 ;
			15'h00000D49 : data <= 8'b00000000 ;
			15'h00000D4A : data <= 8'b00000000 ;
			15'h00000D4B : data <= 8'b00000000 ;
			15'h00000D4C : data <= 8'b00000000 ;
			15'h00000D4D : data <= 8'b00000000 ;
			15'h00000D4E : data <= 8'b00000000 ;
			15'h00000D4F : data <= 8'b00000000 ;
			15'h00000D50 : data <= 8'b00000000 ;
			15'h00000D51 : data <= 8'b00000000 ;
			15'h00000D52 : data <= 8'b00000000 ;
			15'h00000D53 : data <= 8'b00000000 ;
			15'h00000D54 : data <= 8'b00000000 ;
			15'h00000D55 : data <= 8'b00000000 ;
			15'h00000D56 : data <= 8'b00000000 ;
			15'h00000D57 : data <= 8'b00000000 ;
			15'h00000D58 : data <= 8'b00000000 ;
			15'h00000D59 : data <= 8'b00000000 ;
			15'h00000D5A : data <= 8'b00000000 ;
			15'h00000D5B : data <= 8'b00000000 ;
			15'h00000D5C : data <= 8'b00000000 ;
			15'h00000D5D : data <= 8'b00000000 ;
			15'h00000D5E : data <= 8'b00000000 ;
			15'h00000D5F : data <= 8'b00000000 ;
			15'h00000D60 : data <= 8'b00000000 ;
			15'h00000D61 : data <= 8'b00000000 ;
			15'h00000D62 : data <= 8'b00000000 ;
			15'h00000D63 : data <= 8'b00000000 ;
			15'h00000D64 : data <= 8'b00000000 ;
			15'h00000D65 : data <= 8'b00000000 ;
			15'h00000D66 : data <= 8'b00000000 ;
			15'h00000D67 : data <= 8'b00000000 ;
			15'h00000D68 : data <= 8'b00000000 ;
			15'h00000D69 : data <= 8'b00000000 ;
			15'h00000D6A : data <= 8'b00000000 ;
			15'h00000D6B : data <= 8'b00000000 ;
			15'h00000D6C : data <= 8'b00000000 ;
			15'h00000D6D : data <= 8'b00000000 ;
			15'h00000D6E : data <= 8'b00000000 ;
			15'h00000D6F : data <= 8'b00000000 ;
			15'h00000D70 : data <= 8'b00000000 ;
			15'h00000D71 : data <= 8'b00000000 ;
			15'h00000D72 : data <= 8'b00000000 ;
			15'h00000D73 : data <= 8'b00000000 ;
			15'h00000D74 : data <= 8'b00000000 ;
			15'h00000D75 : data <= 8'b00000000 ;
			15'h00000D76 : data <= 8'b00000000 ;
			15'h00000D77 : data <= 8'b00000000 ;
			15'h00000D78 : data <= 8'b00000000 ;
			15'h00000D79 : data <= 8'b00000000 ;
			15'h00000D7A : data <= 8'b00000000 ;
			15'h00000D7B : data <= 8'b00000000 ;
			15'h00000D7C : data <= 8'b00000000 ;
			15'h00000D7D : data <= 8'b00000000 ;
			15'h00000D7E : data <= 8'b00000000 ;
			15'h00000D7F : data <= 8'b00000000 ;
			15'h00000D80 : data <= 8'b00000000 ;
			15'h00000D81 : data <= 8'b00000000 ;
			15'h00000D82 : data <= 8'b00000000 ;
			15'h00000D83 : data <= 8'b00000000 ;
			15'h00000D84 : data <= 8'b00000000 ;
			15'h00000D85 : data <= 8'b00000000 ;
			15'h00000D86 : data <= 8'b00000000 ;
			15'h00000D87 : data <= 8'b00000000 ;
			15'h00000D88 : data <= 8'b00000000 ;
			15'h00000D89 : data <= 8'b00000000 ;
			15'h00000D8A : data <= 8'b00000000 ;
			15'h00000D8B : data <= 8'b00000000 ;
			15'h00000D8C : data <= 8'b00000000 ;
			15'h00000D8D : data <= 8'b00000000 ;
			15'h00000D8E : data <= 8'b00000000 ;
			15'h00000D8F : data <= 8'b00000000 ;
			15'h00000D90 : data <= 8'b00000000 ;
			15'h00000D91 : data <= 8'b00000000 ;
			15'h00000D92 : data <= 8'b00000000 ;
			15'h00000D93 : data <= 8'b00000000 ;
			15'h00000D94 : data <= 8'b00000000 ;
			15'h00000D95 : data <= 8'b00000000 ;
			15'h00000D96 : data <= 8'b00000000 ;
			15'h00000D97 : data <= 8'b00000000 ;
			15'h00000D98 : data <= 8'b00000000 ;
			15'h00000D99 : data <= 8'b00000000 ;
			15'h00000D9A : data <= 8'b00000000 ;
			15'h00000D9B : data <= 8'b00000000 ;
			15'h00000D9C : data <= 8'b00000000 ;
			15'h00000D9D : data <= 8'b00000000 ;
			15'h00000D9E : data <= 8'b00000000 ;
			15'h00000D9F : data <= 8'b00000000 ;
			15'h00000DA0 : data <= 8'b00000000 ;
			15'h00000DA1 : data <= 8'b00000000 ;
			15'h00000DA2 : data <= 8'b00000000 ;
			15'h00000DA3 : data <= 8'b00000000 ;
			15'h00000DA4 : data <= 8'b00000000 ;
			15'h00000DA5 : data <= 8'b00000000 ;
			15'h00000DA6 : data <= 8'b00000000 ;
			15'h00000DA7 : data <= 8'b00000000 ;
			15'h00000DA8 : data <= 8'b00000000 ;
			15'h00000DA9 : data <= 8'b00000000 ;
			15'h00000DAA : data <= 8'b00000000 ;
			15'h00000DAB : data <= 8'b00000000 ;
			15'h00000DAC : data <= 8'b00000000 ;
			15'h00000DAD : data <= 8'b00000000 ;
			15'h00000DAE : data <= 8'b00000000 ;
			15'h00000DAF : data <= 8'b00000000 ;
			15'h00000DB0 : data <= 8'b00000000 ;
			15'h00000DB1 : data <= 8'b00000000 ;
			15'h00000DB2 : data <= 8'b00000000 ;
			15'h00000DB3 : data <= 8'b00000000 ;
			15'h00000DB4 : data <= 8'b00000000 ;
			15'h00000DB5 : data <= 8'b00000000 ;
			15'h00000DB6 : data <= 8'b00000000 ;
			15'h00000DB7 : data <= 8'b00000000 ;
			15'h00000DB8 : data <= 8'b00000000 ;
			15'h00000DB9 : data <= 8'b00000000 ;
			15'h00000DBA : data <= 8'b00000000 ;
			15'h00000DBB : data <= 8'b00000000 ;
			15'h00000DBC : data <= 8'b00000000 ;
			15'h00000DBD : data <= 8'b00000000 ;
			15'h00000DBE : data <= 8'b00000000 ;
			15'h00000DBF : data <= 8'b00000000 ;
			15'h00000DC0 : data <= 8'b00000000 ;
			15'h00000DC1 : data <= 8'b00000000 ;
			15'h00000DC2 : data <= 8'b00000000 ;
			15'h00000DC3 : data <= 8'b00000000 ;
			15'h00000DC4 : data <= 8'b00000000 ;
			15'h00000DC5 : data <= 8'b00000000 ;
			15'h00000DC6 : data <= 8'b00000000 ;
			15'h00000DC7 : data <= 8'b00000000 ;
			15'h00000DC8 : data <= 8'b00000000 ;
			15'h00000DC9 : data <= 8'b00000000 ;
			15'h00000DCA : data <= 8'b00000000 ;
			15'h00000DCB : data <= 8'b00000000 ;
			15'h00000DCC : data <= 8'b00000000 ;
			15'h00000DCD : data <= 8'b00000000 ;
			15'h00000DCE : data <= 8'b00000000 ;
			15'h00000DCF : data <= 8'b00000000 ;
			15'h00000DD0 : data <= 8'b00000000 ;
			15'h00000DD1 : data <= 8'b00000000 ;
			15'h00000DD2 : data <= 8'b00000000 ;
			15'h00000DD3 : data <= 8'b00000000 ;
			15'h00000DD4 : data <= 8'b00000000 ;
			15'h00000DD5 : data <= 8'b00000000 ;
			15'h00000DD6 : data <= 8'b00000000 ;
			15'h00000DD7 : data <= 8'b00000000 ;
			15'h00000DD8 : data <= 8'b00000000 ;
			15'h00000DD9 : data <= 8'b00000000 ;
			15'h00000DDA : data <= 8'b00000000 ;
			15'h00000DDB : data <= 8'b00000000 ;
			15'h00000DDC : data <= 8'b00000000 ;
			15'h00000DDD : data <= 8'b00000000 ;
			15'h00000DDE : data <= 8'b00000000 ;
			15'h00000DDF : data <= 8'b00000000 ;
			15'h00000DE0 : data <= 8'b00000000 ;
			15'h00000DE1 : data <= 8'b00000000 ;
			15'h00000DE2 : data <= 8'b00000000 ;
			15'h00000DE3 : data <= 8'b00000000 ;
			15'h00000DE4 : data <= 8'b00000000 ;
			15'h00000DE5 : data <= 8'b00000000 ;
			15'h00000DE6 : data <= 8'b00000000 ;
			15'h00000DE7 : data <= 8'b00000000 ;
			15'h00000DE8 : data <= 8'b00000000 ;
			15'h00000DE9 : data <= 8'b00000000 ;
			15'h00000DEA : data <= 8'b00000000 ;
			15'h00000DEB : data <= 8'b00000000 ;
			15'h00000DEC : data <= 8'b00000000 ;
			15'h00000DED : data <= 8'b00000000 ;
			15'h00000DEE : data <= 8'b00000000 ;
			15'h00000DEF : data <= 8'b00000000 ;
			15'h00000DF0 : data <= 8'b00000000 ;
			15'h00000DF1 : data <= 8'b00000000 ;
			15'h00000DF2 : data <= 8'b00000000 ;
			15'h00000DF3 : data <= 8'b00000000 ;
			15'h00000DF4 : data <= 8'b00000000 ;
			15'h00000DF5 : data <= 8'b00000000 ;
			15'h00000DF6 : data <= 8'b00000000 ;
			15'h00000DF7 : data <= 8'b00000000 ;
			15'h00000DF8 : data <= 8'b00000000 ;
			15'h00000DF9 : data <= 8'b00000000 ;
			15'h00000DFA : data <= 8'b00000000 ;
			15'h00000DFB : data <= 8'b00000000 ;
			15'h00000DFC : data <= 8'b00000000 ;
			15'h00000DFD : data <= 8'b00000000 ;
			15'h00000DFE : data <= 8'b00000000 ;
			15'h00000DFF : data <= 8'b00000000 ;
			15'h00000E00 : data <= 8'b00000000 ;
			15'h00000E01 : data <= 8'b00000000 ;
			15'h00000E02 : data <= 8'b00000000 ;
			15'h00000E03 : data <= 8'b00000000 ;
			15'h00000E04 : data <= 8'b00000000 ;
			15'h00000E05 : data <= 8'b00000000 ;
			15'h00000E06 : data <= 8'b00000000 ;
			15'h00000E07 : data <= 8'b00000000 ;
			15'h00000E08 : data <= 8'b00000000 ;
			15'h00000E09 : data <= 8'b00000000 ;
			15'h00000E0A : data <= 8'b00000000 ;
			15'h00000E0B : data <= 8'b00000000 ;
			15'h00000E0C : data <= 8'b00000000 ;
			15'h00000E0D : data <= 8'b00000000 ;
			15'h00000E0E : data <= 8'b00000000 ;
			15'h00000E0F : data <= 8'b00000000 ;
			15'h00000E10 : data <= 8'b00000000 ;
			15'h00000E11 : data <= 8'b00000000 ;
			15'h00000E12 : data <= 8'b00000000 ;
			15'h00000E13 : data <= 8'b00000000 ;
			15'h00000E14 : data <= 8'b00000000 ;
			15'h00000E15 : data <= 8'b00000000 ;
			15'h00000E16 : data <= 8'b00000000 ;
			15'h00000E17 : data <= 8'b00000000 ;
			15'h00000E18 : data <= 8'b00000000 ;
			15'h00000E19 : data <= 8'b00000000 ;
			15'h00000E1A : data <= 8'b00000000 ;
			15'h00000E1B : data <= 8'b00000000 ;
			15'h00000E1C : data <= 8'b00000000 ;
			15'h00000E1D : data <= 8'b00000000 ;
			15'h00000E1E : data <= 8'b00000000 ;
			15'h00000E1F : data <= 8'b00000000 ;
			15'h00000E20 : data <= 8'b00000000 ;
			15'h00000E21 : data <= 8'b00000000 ;
			15'h00000E22 : data <= 8'b00000000 ;
			15'h00000E23 : data <= 8'b00000000 ;
			15'h00000E24 : data <= 8'b00000000 ;
			15'h00000E25 : data <= 8'b00000000 ;
			15'h00000E26 : data <= 8'b00000000 ;
			15'h00000E27 : data <= 8'b00000000 ;
			15'h00000E28 : data <= 8'b00000000 ;
			15'h00000E29 : data <= 8'b00000000 ;
			15'h00000E2A : data <= 8'b00000000 ;
			15'h00000E2B : data <= 8'b00000000 ;
			15'h00000E2C : data <= 8'b00000000 ;
			15'h00000E2D : data <= 8'b00000000 ;
			15'h00000E2E : data <= 8'b00000000 ;
			15'h00000E2F : data <= 8'b00000000 ;
			15'h00000E30 : data <= 8'b00000000 ;
			15'h00000E31 : data <= 8'b00000000 ;
			15'h00000E32 : data <= 8'b00000000 ;
			15'h00000E33 : data <= 8'b00000000 ;
			15'h00000E34 : data <= 8'b00000000 ;
			15'h00000E35 : data <= 8'b00000000 ;
			15'h00000E36 : data <= 8'b00000000 ;
			15'h00000E37 : data <= 8'b00000000 ;
			15'h00000E38 : data <= 8'b00000000 ;
			15'h00000E39 : data <= 8'b00000000 ;
			15'h00000E3A : data <= 8'b00000000 ;
			15'h00000E3B : data <= 8'b00000000 ;
			15'h00000E3C : data <= 8'b00000000 ;
			15'h00000E3D : data <= 8'b00000000 ;
			15'h00000E3E : data <= 8'b00000000 ;
			15'h00000E3F : data <= 8'b00000000 ;
			15'h00000E40 : data <= 8'b00000000 ;
			15'h00000E41 : data <= 8'b00000000 ;
			15'h00000E42 : data <= 8'b00000000 ;
			15'h00000E43 : data <= 8'b00000000 ;
			15'h00000E44 : data <= 8'b00000000 ;
			15'h00000E45 : data <= 8'b00000000 ;
			15'h00000E46 : data <= 8'b00000000 ;
			15'h00000E47 : data <= 8'b00000000 ;
			15'h00000E48 : data <= 8'b00000000 ;
			15'h00000E49 : data <= 8'b00000000 ;
			15'h00000E4A : data <= 8'b00000000 ;
			15'h00000E4B : data <= 8'b00000000 ;
			15'h00000E4C : data <= 8'b00000000 ;
			15'h00000E4D : data <= 8'b00000000 ;
			15'h00000E4E : data <= 8'b00000000 ;
			15'h00000E4F : data <= 8'b00000000 ;
			15'h00000E50 : data <= 8'b00000000 ;
			15'h00000E51 : data <= 8'b00000000 ;
			15'h00000E52 : data <= 8'b00000000 ;
			15'h00000E53 : data <= 8'b00000000 ;
			15'h00000E54 : data <= 8'b00000000 ;
			15'h00000E55 : data <= 8'b00000000 ;
			15'h00000E56 : data <= 8'b00000000 ;
			15'h00000E57 : data <= 8'b00000000 ;
			15'h00000E58 : data <= 8'b00000000 ;
			15'h00000E59 : data <= 8'b00000000 ;
			15'h00000E5A : data <= 8'b00000000 ;
			15'h00000E5B : data <= 8'b00000000 ;
			15'h00000E5C : data <= 8'b00000000 ;
			15'h00000E5D : data <= 8'b00000000 ;
			15'h00000E5E : data <= 8'b00000000 ;
			15'h00000E5F : data <= 8'b00000000 ;
			15'h00000E60 : data <= 8'b00000000 ;
			15'h00000E61 : data <= 8'b00000000 ;
			15'h00000E62 : data <= 8'b00000000 ;
			15'h00000E63 : data <= 8'b00000000 ;
			15'h00000E64 : data <= 8'b00000000 ;
			15'h00000E65 : data <= 8'b00000000 ;
			15'h00000E66 : data <= 8'b00000000 ;
			15'h00000E67 : data <= 8'b00000000 ;
			15'h00000E68 : data <= 8'b00000000 ;
			15'h00000E69 : data <= 8'b00000000 ;
			15'h00000E6A : data <= 8'b00000000 ;
			15'h00000E6B : data <= 8'b00000000 ;
			15'h00000E6C : data <= 8'b00000000 ;
			15'h00000E6D : data <= 8'b00000000 ;
			15'h00000E6E : data <= 8'b00000000 ;
			15'h00000E6F : data <= 8'b00000000 ;
			15'h00000E70 : data <= 8'b00000000 ;
			15'h00000E71 : data <= 8'b00000000 ;
			15'h00000E72 : data <= 8'b00000000 ;
			15'h00000E73 : data <= 8'b00000000 ;
			15'h00000E74 : data <= 8'b00000000 ;
			15'h00000E75 : data <= 8'b00000000 ;
			15'h00000E76 : data <= 8'b00000000 ;
			15'h00000E77 : data <= 8'b00000000 ;
			15'h00000E78 : data <= 8'b00000000 ;
			15'h00000E79 : data <= 8'b00000000 ;
			15'h00000E7A : data <= 8'b00000000 ;
			15'h00000E7B : data <= 8'b00000000 ;
			15'h00000E7C : data <= 8'b00000000 ;
			15'h00000E7D : data <= 8'b00000000 ;
			15'h00000E7E : data <= 8'b00000000 ;
			15'h00000E7F : data <= 8'b00000000 ;
			15'h00000E80 : data <= 8'b00000000 ;
			15'h00000E81 : data <= 8'b00000000 ;
			15'h00000E82 : data <= 8'b00000000 ;
			15'h00000E83 : data <= 8'b00000000 ;
			15'h00000E84 : data <= 8'b00000000 ;
			15'h00000E85 : data <= 8'b00000000 ;
			15'h00000E86 : data <= 8'b00000000 ;
			15'h00000E87 : data <= 8'b00000000 ;
			15'h00000E88 : data <= 8'b00000000 ;
			15'h00000E89 : data <= 8'b00000000 ;
			15'h00000E8A : data <= 8'b00000000 ;
			15'h00000E8B : data <= 8'b00000000 ;
			15'h00000E8C : data <= 8'b00000000 ;
			15'h00000E8D : data <= 8'b00000000 ;
			15'h00000E8E : data <= 8'b00000000 ;
			15'h00000E8F : data <= 8'b00000000 ;
			15'h00000E90 : data <= 8'b00000000 ;
			15'h00000E91 : data <= 8'b00000000 ;
			15'h00000E92 : data <= 8'b00000000 ;
			15'h00000E93 : data <= 8'b00000000 ;
			15'h00000E94 : data <= 8'b00000000 ;
			15'h00000E95 : data <= 8'b00000000 ;
			15'h00000E96 : data <= 8'b00000000 ;
			15'h00000E97 : data <= 8'b00000000 ;
			15'h00000E98 : data <= 8'b00000000 ;
			15'h00000E99 : data <= 8'b00000000 ;
			15'h00000E9A : data <= 8'b00000000 ;
			15'h00000E9B : data <= 8'b00000000 ;
			15'h00000E9C : data <= 8'b00000000 ;
			15'h00000E9D : data <= 8'b00000000 ;
			15'h00000E9E : data <= 8'b00000000 ;
			15'h00000E9F : data <= 8'b00000000 ;
			15'h00000EA0 : data <= 8'b00000000 ;
			15'h00000EA1 : data <= 8'b00000000 ;
			15'h00000EA2 : data <= 8'b00000000 ;
			15'h00000EA3 : data <= 8'b00000000 ;
			15'h00000EA4 : data <= 8'b00000000 ;
			15'h00000EA5 : data <= 8'b00000000 ;
			15'h00000EA6 : data <= 8'b00000000 ;
			15'h00000EA7 : data <= 8'b00000000 ;
			15'h00000EA8 : data <= 8'b00000000 ;
			15'h00000EA9 : data <= 8'b00000000 ;
			15'h00000EAA : data <= 8'b00000000 ;
			15'h00000EAB : data <= 8'b00000000 ;
			15'h00000EAC : data <= 8'b00000000 ;
			15'h00000EAD : data <= 8'b00000000 ;
			15'h00000EAE : data <= 8'b00000000 ;
			15'h00000EAF : data <= 8'b00000000 ;
			15'h00000EB0 : data <= 8'b00000000 ;
			15'h00000EB1 : data <= 8'b00000000 ;
			15'h00000EB2 : data <= 8'b00000000 ;
			15'h00000EB3 : data <= 8'b00000000 ;
			15'h00000EB4 : data <= 8'b00000000 ;
			15'h00000EB5 : data <= 8'b00000000 ;
			15'h00000EB6 : data <= 8'b00000000 ;
			15'h00000EB7 : data <= 8'b00000000 ;
			15'h00000EB8 : data <= 8'b00000000 ;
			15'h00000EB9 : data <= 8'b00000000 ;
			15'h00000EBA : data <= 8'b00000000 ;
			15'h00000EBB : data <= 8'b00000000 ;
			15'h00000EBC : data <= 8'b00000000 ;
			15'h00000EBD : data <= 8'b00000000 ;
			15'h00000EBE : data <= 8'b00000000 ;
			15'h00000EBF : data <= 8'b00000000 ;
			15'h00000EC0 : data <= 8'b00000000 ;
			15'h00000EC1 : data <= 8'b00000000 ;
			15'h00000EC2 : data <= 8'b00000000 ;
			15'h00000EC3 : data <= 8'b00000000 ;
			15'h00000EC4 : data <= 8'b00000000 ;
			15'h00000EC5 : data <= 8'b00000000 ;
			15'h00000EC6 : data <= 8'b00000000 ;
			15'h00000EC7 : data <= 8'b00000000 ;
			15'h00000EC8 : data <= 8'b00000000 ;
			15'h00000EC9 : data <= 8'b00000000 ;
			15'h00000ECA : data <= 8'b00000000 ;
			15'h00000ECB : data <= 8'b00000000 ;
			15'h00000ECC : data <= 8'b00000000 ;
			15'h00000ECD : data <= 8'b00000000 ;
			15'h00000ECE : data <= 8'b00000000 ;
			15'h00000ECF : data <= 8'b00000000 ;
			15'h00000ED0 : data <= 8'b00000000 ;
			15'h00000ED1 : data <= 8'b00000000 ;
			15'h00000ED2 : data <= 8'b00000000 ;
			15'h00000ED3 : data <= 8'b00000000 ;
			15'h00000ED4 : data <= 8'b00000000 ;
			15'h00000ED5 : data <= 8'b00000000 ;
			15'h00000ED6 : data <= 8'b00000000 ;
			15'h00000ED7 : data <= 8'b00000000 ;
			15'h00000ED8 : data <= 8'b00000000 ;
			15'h00000ED9 : data <= 8'b00000000 ;
			15'h00000EDA : data <= 8'b00000000 ;
			15'h00000EDB : data <= 8'b00000000 ;
			15'h00000EDC : data <= 8'b00000000 ;
			15'h00000EDD : data <= 8'b00000000 ;
			15'h00000EDE : data <= 8'b00000000 ;
			15'h00000EDF : data <= 8'b00000000 ;
			15'h00000EE0 : data <= 8'b00000000 ;
			15'h00000EE1 : data <= 8'b00000000 ;
			15'h00000EE2 : data <= 8'b00000000 ;
			15'h00000EE3 : data <= 8'b00000000 ;
			15'h00000EE4 : data <= 8'b00000000 ;
			15'h00000EE5 : data <= 8'b00000000 ;
			15'h00000EE6 : data <= 8'b00000000 ;
			15'h00000EE7 : data <= 8'b00000000 ;
			15'h00000EE8 : data <= 8'b00000000 ;
			15'h00000EE9 : data <= 8'b00000000 ;
			15'h00000EEA : data <= 8'b00000000 ;
			15'h00000EEB : data <= 8'b00000000 ;
			15'h00000EEC : data <= 8'b00000000 ;
			15'h00000EED : data <= 8'b00000000 ;
			15'h00000EEE : data <= 8'b00000000 ;
			15'h00000EEF : data <= 8'b00000000 ;
			15'h00000EF0 : data <= 8'b00000000 ;
			15'h00000EF1 : data <= 8'b00000000 ;
			15'h00000EF2 : data <= 8'b00000000 ;
			15'h00000EF3 : data <= 8'b00000000 ;
			15'h00000EF4 : data <= 8'b00000000 ;
			15'h00000EF5 : data <= 8'b00000000 ;
			15'h00000EF6 : data <= 8'b00000000 ;
			15'h00000EF7 : data <= 8'b00000000 ;
			15'h00000EF8 : data <= 8'b00000000 ;
			15'h00000EF9 : data <= 8'b00000000 ;
			15'h00000EFA : data <= 8'b00000000 ;
			15'h00000EFB : data <= 8'b00000000 ;
			15'h00000EFC : data <= 8'b00000000 ;
			15'h00000EFD : data <= 8'b00000000 ;
			15'h00000EFE : data <= 8'b00000000 ;
			15'h00000EFF : data <= 8'b00000000 ;
			15'h00000F00 : data <= 8'b00000000 ;
			15'h00000F01 : data <= 8'b00000000 ;
			15'h00000F02 : data <= 8'b00000000 ;
			15'h00000F03 : data <= 8'b00000000 ;
			15'h00000F04 : data <= 8'b00000000 ;
			15'h00000F05 : data <= 8'b00000000 ;
			15'h00000F06 : data <= 8'b00000000 ;
			15'h00000F07 : data <= 8'b00000000 ;
			15'h00000F08 : data <= 8'b00000000 ;
			15'h00000F09 : data <= 8'b00000000 ;
			15'h00000F0A : data <= 8'b00000000 ;
			15'h00000F0B : data <= 8'b00000000 ;
			15'h00000F0C : data <= 8'b00000000 ;
			15'h00000F0D : data <= 8'b00000000 ;
			15'h00000F0E : data <= 8'b00000000 ;
			15'h00000F0F : data <= 8'b00000000 ;
			15'h00000F10 : data <= 8'b00000000 ;
			15'h00000F11 : data <= 8'b00000000 ;
			15'h00000F12 : data <= 8'b00000000 ;
			15'h00000F13 : data <= 8'b00000000 ;
			15'h00000F14 : data <= 8'b00000000 ;
			15'h00000F15 : data <= 8'b00000000 ;
			15'h00000F16 : data <= 8'b00000000 ;
			15'h00000F17 : data <= 8'b00000000 ;
			15'h00000F18 : data <= 8'b00000000 ;
			15'h00000F19 : data <= 8'b00000000 ;
			15'h00000F1A : data <= 8'b00000000 ;
			15'h00000F1B : data <= 8'b00000000 ;
			15'h00000F1C : data <= 8'b00000000 ;
			15'h00000F1D : data <= 8'b00000000 ;
			15'h00000F1E : data <= 8'b00000000 ;
			15'h00000F1F : data <= 8'b00000000 ;
			15'h00000F20 : data <= 8'b00000000 ;
			15'h00000F21 : data <= 8'b00000000 ;
			15'h00000F22 : data <= 8'b00000000 ;
			15'h00000F23 : data <= 8'b00000000 ;
			15'h00000F24 : data <= 8'b00000000 ;
			15'h00000F25 : data <= 8'b00000000 ;
			15'h00000F26 : data <= 8'b00000000 ;
			15'h00000F27 : data <= 8'b00000000 ;
			15'h00000F28 : data <= 8'b00000000 ;
			15'h00000F29 : data <= 8'b00000000 ;
			15'h00000F2A : data <= 8'b00000000 ;
			15'h00000F2B : data <= 8'b00000000 ;
			15'h00000F2C : data <= 8'b00000000 ;
			15'h00000F2D : data <= 8'b00000000 ;
			15'h00000F2E : data <= 8'b00000000 ;
			15'h00000F2F : data <= 8'b00000000 ;
			15'h00000F30 : data <= 8'b00000000 ;
			15'h00000F31 : data <= 8'b00000000 ;
			15'h00000F32 : data <= 8'b00000000 ;
			15'h00000F33 : data <= 8'b00000000 ;
			15'h00000F34 : data <= 8'b00000000 ;
			15'h00000F35 : data <= 8'b00000000 ;
			15'h00000F36 : data <= 8'b00000000 ;
			15'h00000F37 : data <= 8'b00000000 ;
			15'h00000F38 : data <= 8'b00000000 ;
			15'h00000F39 : data <= 8'b00000000 ;
			15'h00000F3A : data <= 8'b00000000 ;
			15'h00000F3B : data <= 8'b00000000 ;
			15'h00000F3C : data <= 8'b00000000 ;
			15'h00000F3D : data <= 8'b00000000 ;
			15'h00000F3E : data <= 8'b00000000 ;
			15'h00000F3F : data <= 8'b00000000 ;
			15'h00000F40 : data <= 8'b00000000 ;
			15'h00000F41 : data <= 8'b00000000 ;
			15'h00000F42 : data <= 8'b00000000 ;
			15'h00000F43 : data <= 8'b00000000 ;
			15'h00000F44 : data <= 8'b00000000 ;
			15'h00000F45 : data <= 8'b00000000 ;
			15'h00000F46 : data <= 8'b00000000 ;
			15'h00000F47 : data <= 8'b00000000 ;
			15'h00000F48 : data <= 8'b00000000 ;
			15'h00000F49 : data <= 8'b00000000 ;
			15'h00000F4A : data <= 8'b00000000 ;
			15'h00000F4B : data <= 8'b00000000 ;
			15'h00000F4C : data <= 8'b00000000 ;
			15'h00000F4D : data <= 8'b00000000 ;
			15'h00000F4E : data <= 8'b00000000 ;
			15'h00000F4F : data <= 8'b00000000 ;
			15'h00000F50 : data <= 8'b00000000 ;
			15'h00000F51 : data <= 8'b00000000 ;
			15'h00000F52 : data <= 8'b00000000 ;
			15'h00000F53 : data <= 8'b00000000 ;
			15'h00000F54 : data <= 8'b00000000 ;
			15'h00000F55 : data <= 8'b00000000 ;
			15'h00000F56 : data <= 8'b00000000 ;
			15'h00000F57 : data <= 8'b00000000 ;
			15'h00000F58 : data <= 8'b00000000 ;
			15'h00000F59 : data <= 8'b00000000 ;
			15'h00000F5A : data <= 8'b00000000 ;
			15'h00000F5B : data <= 8'b00000000 ;
			15'h00000F5C : data <= 8'b00000000 ;
			15'h00000F5D : data <= 8'b00000000 ;
			15'h00000F5E : data <= 8'b00000000 ;
			15'h00000F5F : data <= 8'b00000000 ;
			15'h00000F60 : data <= 8'b00000000 ;
			15'h00000F61 : data <= 8'b00000000 ;
			15'h00000F62 : data <= 8'b00000000 ;
			15'h00000F63 : data <= 8'b00000000 ;
			15'h00000F64 : data <= 8'b00000000 ;
			15'h00000F65 : data <= 8'b00000000 ;
			15'h00000F66 : data <= 8'b00000000 ;
			15'h00000F67 : data <= 8'b00000000 ;
			15'h00000F68 : data <= 8'b00000000 ;
			15'h00000F69 : data <= 8'b00000000 ;
			15'h00000F6A : data <= 8'b00000000 ;
			15'h00000F6B : data <= 8'b00000000 ;
			15'h00000F6C : data <= 8'b00000000 ;
			15'h00000F6D : data <= 8'b00000000 ;
			15'h00000F6E : data <= 8'b00000000 ;
			15'h00000F6F : data <= 8'b00000000 ;
			15'h00000F70 : data <= 8'b00000000 ;
			15'h00000F71 : data <= 8'b00000000 ;
			15'h00000F72 : data <= 8'b00000000 ;
			15'h00000F73 : data <= 8'b00000000 ;
			15'h00000F74 : data <= 8'b00000000 ;
			15'h00000F75 : data <= 8'b00000000 ;
			15'h00000F76 : data <= 8'b00000000 ;
			15'h00000F77 : data <= 8'b00000000 ;
			15'h00000F78 : data <= 8'b00000000 ;
			15'h00000F79 : data <= 8'b00000000 ;
			15'h00000F7A : data <= 8'b00000000 ;
			15'h00000F7B : data <= 8'b00000000 ;
			15'h00000F7C : data <= 8'b00000000 ;
			15'h00000F7D : data <= 8'b00000000 ;
			15'h00000F7E : data <= 8'b00000000 ;
			15'h00000F7F : data <= 8'b00000000 ;
			15'h00000F80 : data <= 8'b00000000 ;
			15'h00000F81 : data <= 8'b00000000 ;
			15'h00000F82 : data <= 8'b00000000 ;
			15'h00000F83 : data <= 8'b00000000 ;
			15'h00000F84 : data <= 8'b00000000 ;
			15'h00000F85 : data <= 8'b00000000 ;
			15'h00000F86 : data <= 8'b00000000 ;
			15'h00000F87 : data <= 8'b00000000 ;
			15'h00000F88 : data <= 8'b00000000 ;
			15'h00000F89 : data <= 8'b00000000 ;
			15'h00000F8A : data <= 8'b00000000 ;
			15'h00000F8B : data <= 8'b00000000 ;
			15'h00000F8C : data <= 8'b00000000 ;
			15'h00000F8D : data <= 8'b00000000 ;
			15'h00000F8E : data <= 8'b00000000 ;
			15'h00000F8F : data <= 8'b00000000 ;
			15'h00000F90 : data <= 8'b00000000 ;
			15'h00000F91 : data <= 8'b00000000 ;
			15'h00000F92 : data <= 8'b00000000 ;
			15'h00000F93 : data <= 8'b00000000 ;
			15'h00000F94 : data <= 8'b00000000 ;
			15'h00000F95 : data <= 8'b00000000 ;
			15'h00000F96 : data <= 8'b00000000 ;
			15'h00000F97 : data <= 8'b00000000 ;
			15'h00000F98 : data <= 8'b00000000 ;
			15'h00000F99 : data <= 8'b00000000 ;
			15'h00000F9A : data <= 8'b00000000 ;
			15'h00000F9B : data <= 8'b00000000 ;
			15'h00000F9C : data <= 8'b00000000 ;
			15'h00000F9D : data <= 8'b00000000 ;
			15'h00000F9E : data <= 8'b00000000 ;
			15'h00000F9F : data <= 8'b00000000 ;
			15'h00000FA0 : data <= 8'b00000000 ;
			15'h00000FA1 : data <= 8'b00000000 ;
			15'h00000FA2 : data <= 8'b00000000 ;
			15'h00000FA3 : data <= 8'b00000000 ;
			15'h00000FA4 : data <= 8'b00000000 ;
			15'h00000FA5 : data <= 8'b00000000 ;
			15'h00000FA6 : data <= 8'b00000000 ;
			15'h00000FA7 : data <= 8'b00000000 ;
			15'h00000FA8 : data <= 8'b00000000 ;
			15'h00000FA9 : data <= 8'b00000000 ;
			15'h00000FAA : data <= 8'b00000000 ;
			15'h00000FAB : data <= 8'b00000000 ;
			15'h00000FAC : data <= 8'b00000000 ;
			15'h00000FAD : data <= 8'b00000000 ;
			15'h00000FAE : data <= 8'b00000000 ;
			15'h00000FAF : data <= 8'b00000000 ;
			15'h00000FB0 : data <= 8'b00000000 ;
			15'h00000FB1 : data <= 8'b00000000 ;
			15'h00000FB2 : data <= 8'b00000000 ;
			15'h00000FB3 : data <= 8'b00000000 ;
			15'h00000FB4 : data <= 8'b00000000 ;
			15'h00000FB5 : data <= 8'b00000000 ;
			15'h00000FB6 : data <= 8'b00000000 ;
			15'h00000FB7 : data <= 8'b00000000 ;
			15'h00000FB8 : data <= 8'b00000000 ;
			15'h00000FB9 : data <= 8'b00000000 ;
			15'h00000FBA : data <= 8'b00000000 ;
			15'h00000FBB : data <= 8'b00000000 ;
			15'h00000FBC : data <= 8'b00000000 ;
			15'h00000FBD : data <= 8'b00000000 ;
			15'h00000FBE : data <= 8'b00000000 ;
			15'h00000FBF : data <= 8'b00000000 ;
			15'h00000FC0 : data <= 8'b00000000 ;
			15'h00000FC1 : data <= 8'b00000000 ;
			15'h00000FC2 : data <= 8'b00000000 ;
			15'h00000FC3 : data <= 8'b00000000 ;
			15'h00000FC4 : data <= 8'b00000000 ;
			15'h00000FC5 : data <= 8'b00000000 ;
			15'h00000FC6 : data <= 8'b00000000 ;
			15'h00000FC7 : data <= 8'b00000000 ;
			15'h00000FC8 : data <= 8'b00000000 ;
			15'h00000FC9 : data <= 8'b00000000 ;
			15'h00000FCA : data <= 8'b00000000 ;
			15'h00000FCB : data <= 8'b00000000 ;
			15'h00000FCC : data <= 8'b00000000 ;
			15'h00000FCD : data <= 8'b00000000 ;
			15'h00000FCE : data <= 8'b00000000 ;
			15'h00000FCF : data <= 8'b00000000 ;
			15'h00000FD0 : data <= 8'b00000000 ;
			15'h00000FD1 : data <= 8'b00000000 ;
			15'h00000FD2 : data <= 8'b00000000 ;
			15'h00000FD3 : data <= 8'b00000000 ;
			15'h00000FD4 : data <= 8'b00000000 ;
			15'h00000FD5 : data <= 8'b00000000 ;
			15'h00000FD6 : data <= 8'b00000000 ;
			15'h00000FD7 : data <= 8'b00000000 ;
			15'h00000FD8 : data <= 8'b00000000 ;
			15'h00000FD9 : data <= 8'b00000000 ;
			15'h00000FDA : data <= 8'b00000000 ;
			15'h00000FDB : data <= 8'b00000000 ;
			15'h00000FDC : data <= 8'b00000000 ;
			15'h00000FDD : data <= 8'b00000000 ;
			15'h00000FDE : data <= 8'b00000000 ;
			15'h00000FDF : data <= 8'b00000000 ;
			15'h00000FE0 : data <= 8'b00000000 ;
			15'h00000FE1 : data <= 8'b00000000 ;
			15'h00000FE2 : data <= 8'b00000000 ;
			15'h00000FE3 : data <= 8'b00000000 ;
			15'h00000FE4 : data <= 8'b00000000 ;
			15'h00000FE5 : data <= 8'b00000000 ;
			15'h00000FE6 : data <= 8'b00000000 ;
			15'h00000FE7 : data <= 8'b00000000 ;
			15'h00000FE8 : data <= 8'b00000000 ;
			15'h00000FE9 : data <= 8'b00000000 ;
			15'h00000FEA : data <= 8'b00000000 ;
			15'h00000FEB : data <= 8'b00000000 ;
			15'h00000FEC : data <= 8'b00000000 ;
			15'h00000FED : data <= 8'b00000000 ;
			15'h00000FEE : data <= 8'b00000000 ;
			15'h00000FEF : data <= 8'b00000000 ;
			15'h00000FF0 : data <= 8'b00000000 ;
			15'h00000FF1 : data <= 8'b00000000 ;
			15'h00000FF2 : data <= 8'b00000000 ;
			15'h00000FF3 : data <= 8'b00000000 ;
			15'h00000FF4 : data <= 8'b00000000 ;
			15'h00000FF5 : data <= 8'b00000000 ;
			15'h00000FF6 : data <= 8'b00000000 ;
			15'h00000FF7 : data <= 8'b00000000 ;
			15'h00000FF8 : data <= 8'b00000000 ;
			15'h00000FF9 : data <= 8'b00000000 ;
			15'h00000FFA : data <= 8'b00000000 ;
			15'h00000FFB : data <= 8'b00000000 ;
			15'h00000FFC : data <= 8'b00000000 ;
			15'h00000FFD : data <= 8'b00000000 ;
			15'h00000FFE : data <= 8'b00000000 ;
			15'h00000FFF : data <= 8'b00000000 ;
			15'h00001000 : data <= 8'b00000000 ;
			15'h00001001 : data <= 8'b00000000 ;
			15'h00001002 : data <= 8'b00000000 ;
			15'h00001003 : data <= 8'b00000000 ;
			15'h00001004 : data <= 8'b00000000 ;
			15'h00001005 : data <= 8'b00000000 ;
			15'h00001006 : data <= 8'b00000000 ;
			15'h00001007 : data <= 8'b00000000 ;
			15'h00001008 : data <= 8'b00000000 ;
			15'h00001009 : data <= 8'b00000000 ;
			15'h0000100A : data <= 8'b00000000 ;
			15'h0000100B : data <= 8'b00000000 ;
			15'h0000100C : data <= 8'b00000000 ;
			15'h0000100D : data <= 8'b00000000 ;
			15'h0000100E : data <= 8'b00000000 ;
			15'h0000100F : data <= 8'b00000000 ;
			15'h00001010 : data <= 8'b00000000 ;
			15'h00001011 : data <= 8'b00000000 ;
			15'h00001012 : data <= 8'b00000000 ;
			15'h00001013 : data <= 8'b00000000 ;
			15'h00001014 : data <= 8'b00000000 ;
			15'h00001015 : data <= 8'b00000000 ;
			15'h00001016 : data <= 8'b00000000 ;
			15'h00001017 : data <= 8'b00000000 ;
			15'h00001018 : data <= 8'b00000000 ;
			15'h00001019 : data <= 8'b00000000 ;
			15'h0000101A : data <= 8'b00000000 ;
			15'h0000101B : data <= 8'b00000000 ;
			15'h0000101C : data <= 8'b00000000 ;
			15'h0000101D : data <= 8'b00000000 ;
			15'h0000101E : data <= 8'b00000000 ;
			15'h0000101F : data <= 8'b00000000 ;
			15'h00001020 : data <= 8'b00000000 ;
			15'h00001021 : data <= 8'b00000000 ;
			15'h00001022 : data <= 8'b00000000 ;
			15'h00001023 : data <= 8'b00000000 ;
			15'h00001024 : data <= 8'b00000000 ;
			15'h00001025 : data <= 8'b00000000 ;
			15'h00001026 : data <= 8'b00000000 ;
			15'h00001027 : data <= 8'b00000000 ;
			15'h00001028 : data <= 8'b00000000 ;
			15'h00001029 : data <= 8'b00000000 ;
			15'h0000102A : data <= 8'b00000000 ;
			15'h0000102B : data <= 8'b00000000 ;
			15'h0000102C : data <= 8'b00000000 ;
			15'h0000102D : data <= 8'b00000000 ;
			15'h0000102E : data <= 8'b00000000 ;
			15'h0000102F : data <= 8'b00000000 ;
			15'h00001030 : data <= 8'b00000000 ;
			15'h00001031 : data <= 8'b00000000 ;
			15'h00001032 : data <= 8'b00000000 ;
			15'h00001033 : data <= 8'b00000000 ;
			15'h00001034 : data <= 8'b00000000 ;
			15'h00001035 : data <= 8'b00000000 ;
			15'h00001036 : data <= 8'b00000000 ;
			15'h00001037 : data <= 8'b00000000 ;
			15'h00001038 : data <= 8'b00000000 ;
			15'h00001039 : data <= 8'b00000000 ;
			15'h0000103A : data <= 8'b00000000 ;
			15'h0000103B : data <= 8'b00000000 ;
			15'h0000103C : data <= 8'b00000000 ;
			15'h0000103D : data <= 8'b00000000 ;
			15'h0000103E : data <= 8'b00000000 ;
			15'h0000103F : data <= 8'b00000000 ;
			15'h00001040 : data <= 8'b00000000 ;
			15'h00001041 : data <= 8'b00000000 ;
			15'h00001042 : data <= 8'b00000000 ;
			15'h00001043 : data <= 8'b00000000 ;
			15'h00001044 : data <= 8'b00000000 ;
			15'h00001045 : data <= 8'b00000000 ;
			15'h00001046 : data <= 8'b00000000 ;
			15'h00001047 : data <= 8'b00000000 ;
			15'h00001048 : data <= 8'b00000000 ;
			15'h00001049 : data <= 8'b00000000 ;
			15'h0000104A : data <= 8'b00000000 ;
			15'h0000104B : data <= 8'b00000000 ;
			15'h0000104C : data <= 8'b00000000 ;
			15'h0000104D : data <= 8'b00000000 ;
			15'h0000104E : data <= 8'b00000000 ;
			15'h0000104F : data <= 8'b00000000 ;
			15'h00001050 : data <= 8'b00000000 ;
			15'h00001051 : data <= 8'b00000000 ;
			15'h00001052 : data <= 8'b00000000 ;
			15'h00001053 : data <= 8'b00000000 ;
			15'h00001054 : data <= 8'b00000000 ;
			15'h00001055 : data <= 8'b00000000 ;
			15'h00001056 : data <= 8'b00000000 ;
			15'h00001057 : data <= 8'b00000000 ;
			15'h00001058 : data <= 8'b00000000 ;
			15'h00001059 : data <= 8'b00000000 ;
			15'h0000105A : data <= 8'b00000000 ;
			15'h0000105B : data <= 8'b00000000 ;
			15'h0000105C : data <= 8'b00000000 ;
			15'h0000105D : data <= 8'b00000000 ;
			15'h0000105E : data <= 8'b00000000 ;
			15'h0000105F : data <= 8'b00000000 ;
			15'h00001060 : data <= 8'b00000000 ;
			15'h00001061 : data <= 8'b00000000 ;
			15'h00001062 : data <= 8'b00000000 ;
			15'h00001063 : data <= 8'b00000000 ;
			15'h00001064 : data <= 8'b00000000 ;
			15'h00001065 : data <= 8'b00000000 ;
			15'h00001066 : data <= 8'b00000000 ;
			15'h00001067 : data <= 8'b00000000 ;
			15'h00001068 : data <= 8'b00000000 ;
			15'h00001069 : data <= 8'b00000000 ;
			15'h0000106A : data <= 8'b00000000 ;
			15'h0000106B : data <= 8'b00000000 ;
			15'h0000106C : data <= 8'b00000000 ;
			15'h0000106D : data <= 8'b00000000 ;
			15'h0000106E : data <= 8'b00000000 ;
			15'h0000106F : data <= 8'b00000000 ;
			15'h00001070 : data <= 8'b00000000 ;
			15'h00001071 : data <= 8'b00000000 ;
			15'h00001072 : data <= 8'b00000000 ;
			15'h00001073 : data <= 8'b00000000 ;
			15'h00001074 : data <= 8'b00000000 ;
			15'h00001075 : data <= 8'b00000000 ;
			15'h00001076 : data <= 8'b00000000 ;
			15'h00001077 : data <= 8'b00000000 ;
			15'h00001078 : data <= 8'b00000000 ;
			15'h00001079 : data <= 8'b00000000 ;
			15'h0000107A : data <= 8'b00000000 ;
			15'h0000107B : data <= 8'b00000000 ;
			15'h0000107C : data <= 8'b00000000 ;
			15'h0000107D : data <= 8'b00000000 ;
			15'h0000107E : data <= 8'b00000000 ;
			15'h0000107F : data <= 8'b00000000 ;
			15'h00001080 : data <= 8'b00000000 ;
			15'h00001081 : data <= 8'b00000000 ;
			15'h00001082 : data <= 8'b00000000 ;
			15'h00001083 : data <= 8'b00000000 ;
			15'h00001084 : data <= 8'b00000000 ;
			15'h00001085 : data <= 8'b00000000 ;
			15'h00001086 : data <= 8'b00000000 ;
			15'h00001087 : data <= 8'b00000000 ;
			15'h00001088 : data <= 8'b00000000 ;
			15'h00001089 : data <= 8'b00000000 ;
			15'h0000108A : data <= 8'b00000000 ;
			15'h0000108B : data <= 8'b00000000 ;
			15'h0000108C : data <= 8'b00000000 ;
			15'h0000108D : data <= 8'b00000000 ;
			15'h0000108E : data <= 8'b00000000 ;
			15'h0000108F : data <= 8'b00000000 ;
			15'h00001090 : data <= 8'b00000000 ;
			15'h00001091 : data <= 8'b00000000 ;
			15'h00001092 : data <= 8'b00000000 ;
			15'h00001093 : data <= 8'b00000000 ;
			15'h00001094 : data <= 8'b00000000 ;
			15'h00001095 : data <= 8'b00000000 ;
			15'h00001096 : data <= 8'b00000000 ;
			15'h00001097 : data <= 8'b00000000 ;
			15'h00001098 : data <= 8'b00000000 ;
			15'h00001099 : data <= 8'b00000000 ;
			15'h0000109A : data <= 8'b00000000 ;
			15'h0000109B : data <= 8'b00000000 ;
			15'h0000109C : data <= 8'b00000000 ;
			15'h0000109D : data <= 8'b00000000 ;
			15'h0000109E : data <= 8'b00000000 ;
			15'h0000109F : data <= 8'b00000000 ;
			15'h000010A0 : data <= 8'b00000000 ;
			15'h000010A1 : data <= 8'b00000000 ;
			15'h000010A2 : data <= 8'b00000000 ;
			15'h000010A3 : data <= 8'b00000000 ;
			15'h000010A4 : data <= 8'b00000000 ;
			15'h000010A5 : data <= 8'b00000000 ;
			15'h000010A6 : data <= 8'b00000000 ;
			15'h000010A7 : data <= 8'b00000000 ;
			15'h000010A8 : data <= 8'b00000000 ;
			15'h000010A9 : data <= 8'b00000000 ;
			15'h000010AA : data <= 8'b00000000 ;
			15'h000010AB : data <= 8'b00000000 ;
			15'h000010AC : data <= 8'b00000000 ;
			15'h000010AD : data <= 8'b00000000 ;
			15'h000010AE : data <= 8'b00000000 ;
			15'h000010AF : data <= 8'b00000000 ;
			15'h000010B0 : data <= 8'b00000000 ;
			15'h000010B1 : data <= 8'b00000000 ;
			15'h000010B2 : data <= 8'b00000000 ;
			15'h000010B3 : data <= 8'b00000000 ;
			15'h000010B4 : data <= 8'b00000000 ;
			15'h000010B5 : data <= 8'b00000000 ;
			15'h000010B6 : data <= 8'b00000000 ;
			15'h000010B7 : data <= 8'b00000000 ;
			15'h000010B8 : data <= 8'b00000000 ;
			15'h000010B9 : data <= 8'b00000000 ;
			15'h000010BA : data <= 8'b00000000 ;
			15'h000010BB : data <= 8'b00000000 ;
			15'h000010BC : data <= 8'b00000000 ;
			15'h000010BD : data <= 8'b00000000 ;
			15'h000010BE : data <= 8'b00000000 ;
			15'h000010BF : data <= 8'b00000000 ;
			15'h000010C0 : data <= 8'b00000000 ;
			15'h000010C1 : data <= 8'b00000000 ;
			15'h000010C2 : data <= 8'b00000000 ;
			15'h000010C3 : data <= 8'b00000000 ;
			15'h000010C4 : data <= 8'b00000000 ;
			15'h000010C5 : data <= 8'b00000000 ;
			15'h000010C6 : data <= 8'b00000000 ;
			15'h000010C7 : data <= 8'b00000000 ;
			15'h000010C8 : data <= 8'b00000000 ;
			15'h000010C9 : data <= 8'b00000000 ;
			15'h000010CA : data <= 8'b00000000 ;
			15'h000010CB : data <= 8'b00000000 ;
			15'h000010CC : data <= 8'b00000000 ;
			15'h000010CD : data <= 8'b00000000 ;
			15'h000010CE : data <= 8'b00000000 ;
			15'h000010CF : data <= 8'b00000000 ;
			15'h000010D0 : data <= 8'b00000000 ;
			15'h000010D1 : data <= 8'b00000000 ;
			15'h000010D2 : data <= 8'b00000000 ;
			15'h000010D3 : data <= 8'b00000000 ;
			15'h000010D4 : data <= 8'b00000000 ;
			15'h000010D5 : data <= 8'b00000000 ;
			15'h000010D6 : data <= 8'b00000000 ;
			15'h000010D7 : data <= 8'b00000000 ;
			15'h000010D8 : data <= 8'b00000000 ;
			15'h000010D9 : data <= 8'b00000000 ;
			15'h000010DA : data <= 8'b00000000 ;
			15'h000010DB : data <= 8'b00000000 ;
			15'h000010DC : data <= 8'b00000000 ;
			15'h000010DD : data <= 8'b00000000 ;
			15'h000010DE : data <= 8'b00000000 ;
			15'h000010DF : data <= 8'b00000000 ;
			15'h000010E0 : data <= 8'b00000000 ;
			15'h000010E1 : data <= 8'b00000000 ;
			15'h000010E2 : data <= 8'b00000000 ;
			15'h000010E3 : data <= 8'b00000000 ;
			15'h000010E4 : data <= 8'b00000000 ;
			15'h000010E5 : data <= 8'b00000000 ;
			15'h000010E6 : data <= 8'b00000000 ;
			15'h000010E7 : data <= 8'b00000000 ;
			15'h000010E8 : data <= 8'b00000000 ;
			15'h000010E9 : data <= 8'b00000000 ;
			15'h000010EA : data <= 8'b00000000 ;
			15'h000010EB : data <= 8'b00000000 ;
			15'h000010EC : data <= 8'b00000000 ;
			15'h000010ED : data <= 8'b00000000 ;
			15'h000010EE : data <= 8'b00000000 ;
			15'h000010EF : data <= 8'b00000000 ;
			15'h000010F0 : data <= 8'b00000000 ;
			15'h000010F1 : data <= 8'b00000000 ;
			15'h000010F2 : data <= 8'b00000000 ;
			15'h000010F3 : data <= 8'b00000000 ;
			15'h000010F4 : data <= 8'b00000000 ;
			15'h000010F5 : data <= 8'b00000000 ;
			15'h000010F6 : data <= 8'b00000000 ;
			15'h000010F7 : data <= 8'b00000000 ;
			15'h000010F8 : data <= 8'b00000000 ;
			15'h000010F9 : data <= 8'b00000000 ;
			15'h000010FA : data <= 8'b00000000 ;
			15'h000010FB : data <= 8'b00000000 ;
			15'h000010FC : data <= 8'b00000000 ;
			15'h000010FD : data <= 8'b00000000 ;
			15'h000010FE : data <= 8'b00000000 ;
			15'h000010FF : data <= 8'b00000000 ;
			15'h00001100 : data <= 8'b00000000 ;
			15'h00001101 : data <= 8'b00000000 ;
			15'h00001102 : data <= 8'b00000000 ;
			15'h00001103 : data <= 8'b00000000 ;
			15'h00001104 : data <= 8'b00000000 ;
			15'h00001105 : data <= 8'b00000000 ;
			15'h00001106 : data <= 8'b00000000 ;
			15'h00001107 : data <= 8'b00000000 ;
			15'h00001108 : data <= 8'b00000000 ;
			15'h00001109 : data <= 8'b00000000 ;
			15'h0000110A : data <= 8'b00000000 ;
			15'h0000110B : data <= 8'b00000000 ;
			15'h0000110C : data <= 8'b00000000 ;
			15'h0000110D : data <= 8'b00000000 ;
			15'h0000110E : data <= 8'b00000000 ;
			15'h0000110F : data <= 8'b00000000 ;
			15'h00001110 : data <= 8'b00000000 ;
			15'h00001111 : data <= 8'b00000000 ;
			15'h00001112 : data <= 8'b00000000 ;
			15'h00001113 : data <= 8'b00000000 ;
			15'h00001114 : data <= 8'b00000000 ;
			15'h00001115 : data <= 8'b00000000 ;
			15'h00001116 : data <= 8'b00000000 ;
			15'h00001117 : data <= 8'b00000000 ;
			15'h00001118 : data <= 8'b00000000 ;
			15'h00001119 : data <= 8'b00000000 ;
			15'h0000111A : data <= 8'b00000000 ;
			15'h0000111B : data <= 8'b00000000 ;
			15'h0000111C : data <= 8'b00000000 ;
			15'h0000111D : data <= 8'b00000000 ;
			15'h0000111E : data <= 8'b00000000 ;
			15'h0000111F : data <= 8'b00000000 ;
			15'h00001120 : data <= 8'b00000000 ;
			15'h00001121 : data <= 8'b00000000 ;
			15'h00001122 : data <= 8'b00000000 ;
			15'h00001123 : data <= 8'b00000000 ;
			15'h00001124 : data <= 8'b00000000 ;
			15'h00001125 : data <= 8'b00000000 ;
			15'h00001126 : data <= 8'b00000000 ;
			15'h00001127 : data <= 8'b00000000 ;
			15'h00001128 : data <= 8'b00000000 ;
			15'h00001129 : data <= 8'b00000000 ;
			15'h0000112A : data <= 8'b00000000 ;
			15'h0000112B : data <= 8'b00000000 ;
			15'h0000112C : data <= 8'b00000000 ;
			15'h0000112D : data <= 8'b00000000 ;
			15'h0000112E : data <= 8'b00000000 ;
			15'h0000112F : data <= 8'b00000000 ;
			15'h00001130 : data <= 8'b00000000 ;
			15'h00001131 : data <= 8'b00000000 ;
			15'h00001132 : data <= 8'b00000000 ;
			15'h00001133 : data <= 8'b00000000 ;
			15'h00001134 : data <= 8'b00000000 ;
			15'h00001135 : data <= 8'b00000000 ;
			15'h00001136 : data <= 8'b00000000 ;
			15'h00001137 : data <= 8'b00000000 ;
			15'h00001138 : data <= 8'b00000000 ;
			15'h00001139 : data <= 8'b00000000 ;
			15'h0000113A : data <= 8'b00000000 ;
			15'h0000113B : data <= 8'b00000000 ;
			15'h0000113C : data <= 8'b00000000 ;
			15'h0000113D : data <= 8'b00000000 ;
			15'h0000113E : data <= 8'b00000000 ;
			15'h0000113F : data <= 8'b00000000 ;
			15'h00001140 : data <= 8'b00000000 ;
			15'h00001141 : data <= 8'b00000000 ;
			15'h00001142 : data <= 8'b00000000 ;
			15'h00001143 : data <= 8'b00000000 ;
			15'h00001144 : data <= 8'b00000000 ;
			15'h00001145 : data <= 8'b00000000 ;
			15'h00001146 : data <= 8'b00000000 ;
			15'h00001147 : data <= 8'b00000000 ;
			15'h00001148 : data <= 8'b00000000 ;
			15'h00001149 : data <= 8'b00000000 ;
			15'h0000114A : data <= 8'b00000000 ;
			15'h0000114B : data <= 8'b00000000 ;
			15'h0000114C : data <= 8'b00000000 ;
			15'h0000114D : data <= 8'b00000000 ;
			15'h0000114E : data <= 8'b00000000 ;
			15'h0000114F : data <= 8'b00000000 ;
			15'h00001150 : data <= 8'b00000000 ;
			15'h00001151 : data <= 8'b00000000 ;
			15'h00001152 : data <= 8'b00000000 ;
			15'h00001153 : data <= 8'b00000000 ;
			15'h00001154 : data <= 8'b00000000 ;
			15'h00001155 : data <= 8'b00000000 ;
			15'h00001156 : data <= 8'b00000000 ;
			15'h00001157 : data <= 8'b00000000 ;
			15'h00001158 : data <= 8'b00000000 ;
			15'h00001159 : data <= 8'b00000000 ;
			15'h0000115A : data <= 8'b00000000 ;
			15'h0000115B : data <= 8'b00000000 ;
			15'h0000115C : data <= 8'b00000000 ;
			15'h0000115D : data <= 8'b00000000 ;
			15'h0000115E : data <= 8'b00000000 ;
			15'h0000115F : data <= 8'b00000000 ;
			15'h00001160 : data <= 8'b00000000 ;
			15'h00001161 : data <= 8'b00000000 ;
			15'h00001162 : data <= 8'b00000000 ;
			15'h00001163 : data <= 8'b00000000 ;
			15'h00001164 : data <= 8'b00000000 ;
			15'h00001165 : data <= 8'b00000000 ;
			15'h00001166 : data <= 8'b00000000 ;
			15'h00001167 : data <= 8'b00000000 ;
			15'h00001168 : data <= 8'b00000000 ;
			15'h00001169 : data <= 8'b00000000 ;
			15'h0000116A : data <= 8'b00000000 ;
			15'h0000116B : data <= 8'b00000000 ;
			15'h0000116C : data <= 8'b00000000 ;
			15'h0000116D : data <= 8'b00000000 ;
			15'h0000116E : data <= 8'b00000000 ;
			15'h0000116F : data <= 8'b00000000 ;
			15'h00001170 : data <= 8'b00000000 ;
			15'h00001171 : data <= 8'b00000000 ;
			15'h00001172 : data <= 8'b00000000 ;
			15'h00001173 : data <= 8'b00000000 ;
			15'h00001174 : data <= 8'b00000000 ;
			15'h00001175 : data <= 8'b00000000 ;
			15'h00001176 : data <= 8'b00000000 ;
			15'h00001177 : data <= 8'b00000000 ;
			15'h00001178 : data <= 8'b00000000 ;
			15'h00001179 : data <= 8'b00000000 ;
			15'h0000117A : data <= 8'b00000000 ;
			15'h0000117B : data <= 8'b00000000 ;
			15'h0000117C : data <= 8'b00000000 ;
			15'h0000117D : data <= 8'b00000000 ;
			15'h0000117E : data <= 8'b00000000 ;
			15'h0000117F : data <= 8'b00000000 ;
			15'h00001180 : data <= 8'b00000000 ;
			15'h00001181 : data <= 8'b00000000 ;
			15'h00001182 : data <= 8'b00000000 ;
			15'h00001183 : data <= 8'b00000000 ;
			15'h00001184 : data <= 8'b00000000 ;
			15'h00001185 : data <= 8'b00000000 ;
			15'h00001186 : data <= 8'b00000000 ;
			15'h00001187 : data <= 8'b00000000 ;
			15'h00001188 : data <= 8'b00000000 ;
			15'h00001189 : data <= 8'b00000000 ;
			15'h0000118A : data <= 8'b00000000 ;
			15'h0000118B : data <= 8'b00000000 ;
			15'h0000118C : data <= 8'b00000000 ;
			15'h0000118D : data <= 8'b00000000 ;
			15'h0000118E : data <= 8'b00000000 ;
			15'h0000118F : data <= 8'b00000000 ;
			15'h00001190 : data <= 8'b00000000 ;
			15'h00001191 : data <= 8'b00000000 ;
			15'h00001192 : data <= 8'b00000000 ;
			15'h00001193 : data <= 8'b00000000 ;
			15'h00001194 : data <= 8'b00000000 ;
			15'h00001195 : data <= 8'b00000000 ;
			15'h00001196 : data <= 8'b00000000 ;
			15'h00001197 : data <= 8'b00000000 ;
			15'h00001198 : data <= 8'b00000000 ;
			15'h00001199 : data <= 8'b00000000 ;
			15'h0000119A : data <= 8'b00000000 ;
			15'h0000119B : data <= 8'b00000000 ;
			15'h0000119C : data <= 8'b00000000 ;
			15'h0000119D : data <= 8'b00000000 ;
			15'h0000119E : data <= 8'b00000000 ;
			15'h0000119F : data <= 8'b00000000 ;
			15'h000011A0 : data <= 8'b00000000 ;
			15'h000011A1 : data <= 8'b00000000 ;
			15'h000011A2 : data <= 8'b00000000 ;
			15'h000011A3 : data <= 8'b00000000 ;
			15'h000011A4 : data <= 8'b00000000 ;
			15'h000011A5 : data <= 8'b00000000 ;
			15'h000011A6 : data <= 8'b00000000 ;
			15'h000011A7 : data <= 8'b00000000 ;
			15'h000011A8 : data <= 8'b00000000 ;
			15'h000011A9 : data <= 8'b00000000 ;
			15'h000011AA : data <= 8'b00000000 ;
			15'h000011AB : data <= 8'b00000000 ;
			15'h000011AC : data <= 8'b00000000 ;
			15'h000011AD : data <= 8'b00000000 ;
			15'h000011AE : data <= 8'b00000000 ;
			15'h000011AF : data <= 8'b00000000 ;
			15'h000011B0 : data <= 8'b00000000 ;
			15'h000011B1 : data <= 8'b00000000 ;
			15'h000011B2 : data <= 8'b00000000 ;
			15'h000011B3 : data <= 8'b00000000 ;
			15'h000011B4 : data <= 8'b00000000 ;
			15'h000011B5 : data <= 8'b00000000 ;
			15'h000011B6 : data <= 8'b00000000 ;
			15'h000011B7 : data <= 8'b00000000 ;
			15'h000011B8 : data <= 8'b00000000 ;
			15'h000011B9 : data <= 8'b00000000 ;
			15'h000011BA : data <= 8'b00000000 ;
			15'h000011BB : data <= 8'b00000000 ;
			15'h000011BC : data <= 8'b00000000 ;
			15'h000011BD : data <= 8'b00000000 ;
			15'h000011BE : data <= 8'b00000000 ;
			15'h000011BF : data <= 8'b00000000 ;
			15'h000011C0 : data <= 8'b00000000 ;
			15'h000011C1 : data <= 8'b00000000 ;
			15'h000011C2 : data <= 8'b00000000 ;
			15'h000011C3 : data <= 8'b00000000 ;
			15'h000011C4 : data <= 8'b00000000 ;
			15'h000011C5 : data <= 8'b00000000 ;
			15'h000011C6 : data <= 8'b00000000 ;
			15'h000011C7 : data <= 8'b00000000 ;
			15'h000011C8 : data <= 8'b00000000 ;
			15'h000011C9 : data <= 8'b00000000 ;
			15'h000011CA : data <= 8'b00000000 ;
			15'h000011CB : data <= 8'b00000000 ;
			15'h000011CC : data <= 8'b00000000 ;
			15'h000011CD : data <= 8'b00000000 ;
			15'h000011CE : data <= 8'b00000000 ;
			15'h000011CF : data <= 8'b00000000 ;
			15'h000011D0 : data <= 8'b00000000 ;
			15'h000011D1 : data <= 8'b00000000 ;
			15'h000011D2 : data <= 8'b00000000 ;
			15'h000011D3 : data <= 8'b00000000 ;
			15'h000011D4 : data <= 8'b00000000 ;
			15'h000011D5 : data <= 8'b00000000 ;
			15'h000011D6 : data <= 8'b00000000 ;
			15'h000011D7 : data <= 8'b00000000 ;
			15'h000011D8 : data <= 8'b00000000 ;
			15'h000011D9 : data <= 8'b00000000 ;
			15'h000011DA : data <= 8'b00000000 ;
			15'h000011DB : data <= 8'b00000000 ;
			15'h000011DC : data <= 8'b00000000 ;
			15'h000011DD : data <= 8'b00000000 ;
			15'h000011DE : data <= 8'b00000000 ;
			15'h000011DF : data <= 8'b00000000 ;
			15'h000011E0 : data <= 8'b00000000 ;
			15'h000011E1 : data <= 8'b00000000 ;
			15'h000011E2 : data <= 8'b00000000 ;
			15'h000011E3 : data <= 8'b00000000 ;
			15'h000011E4 : data <= 8'b00000000 ;
			15'h000011E5 : data <= 8'b00000000 ;
			15'h000011E6 : data <= 8'b00000000 ;
			15'h000011E7 : data <= 8'b00000000 ;
			15'h000011E8 : data <= 8'b00000000 ;
			15'h000011E9 : data <= 8'b00000000 ;
			15'h000011EA : data <= 8'b00000000 ;
			15'h000011EB : data <= 8'b00000000 ;
			15'h000011EC : data <= 8'b00000000 ;
			15'h000011ED : data <= 8'b00000000 ;
			15'h000011EE : data <= 8'b00000000 ;
			15'h000011EF : data <= 8'b00000000 ;
			15'h000011F0 : data <= 8'b00000000 ;
			15'h000011F1 : data <= 8'b00000000 ;
			15'h000011F2 : data <= 8'b00000000 ;
			15'h000011F3 : data <= 8'b00000000 ;
			15'h000011F4 : data <= 8'b00000000 ;
			15'h000011F5 : data <= 8'b00000000 ;
			15'h000011F6 : data <= 8'b00000000 ;
			15'h000011F7 : data <= 8'b00000000 ;
			15'h000011F8 : data <= 8'b00000000 ;
			15'h000011F9 : data <= 8'b00000000 ;
			15'h000011FA : data <= 8'b00000000 ;
			15'h000011FB : data <= 8'b00000000 ;
			15'h000011FC : data <= 8'b00000000 ;
			15'h000011FD : data <= 8'b00000000 ;
			15'h000011FE : data <= 8'b00000000 ;
			15'h000011FF : data <= 8'b00000000 ;
			15'h00001200 : data <= 8'b00000000 ;
			15'h00001201 : data <= 8'b00000000 ;
			15'h00001202 : data <= 8'b00000000 ;
			15'h00001203 : data <= 8'b00000000 ;
			15'h00001204 : data <= 8'b00000000 ;
			15'h00001205 : data <= 8'b00000000 ;
			15'h00001206 : data <= 8'b00000000 ;
			15'h00001207 : data <= 8'b00000000 ;
			15'h00001208 : data <= 8'b00000000 ;
			15'h00001209 : data <= 8'b00000000 ;
			15'h0000120A : data <= 8'b00000000 ;
			15'h0000120B : data <= 8'b00000000 ;
			15'h0000120C : data <= 8'b00000000 ;
			15'h0000120D : data <= 8'b00000000 ;
			15'h0000120E : data <= 8'b00000000 ;
			15'h0000120F : data <= 8'b00000000 ;
			15'h00001210 : data <= 8'b00000000 ;
			15'h00001211 : data <= 8'b00000000 ;
			15'h00001212 : data <= 8'b00000000 ;
			15'h00001213 : data <= 8'b00000000 ;
			15'h00001214 : data <= 8'b00000000 ;
			15'h00001215 : data <= 8'b00000000 ;
			15'h00001216 : data <= 8'b00000000 ;
			15'h00001217 : data <= 8'b00000000 ;
			15'h00001218 : data <= 8'b00000000 ;
			15'h00001219 : data <= 8'b00000000 ;
			15'h0000121A : data <= 8'b00000000 ;
			15'h0000121B : data <= 8'b00000000 ;
			15'h0000121C : data <= 8'b00000000 ;
			15'h0000121D : data <= 8'b00000000 ;
			15'h0000121E : data <= 8'b00000000 ;
			15'h0000121F : data <= 8'b00000000 ;
			15'h00001220 : data <= 8'b00000000 ;
			15'h00001221 : data <= 8'b00000000 ;
			15'h00001222 : data <= 8'b00000000 ;
			15'h00001223 : data <= 8'b00000000 ;
			15'h00001224 : data <= 8'b00000000 ;
			15'h00001225 : data <= 8'b00000000 ;
			15'h00001226 : data <= 8'b00000000 ;
			15'h00001227 : data <= 8'b00000000 ;
			15'h00001228 : data <= 8'b00000000 ;
			15'h00001229 : data <= 8'b00000000 ;
			15'h0000122A : data <= 8'b00000000 ;
			15'h0000122B : data <= 8'b00000000 ;
			15'h0000122C : data <= 8'b00000000 ;
			15'h0000122D : data <= 8'b00000000 ;
			15'h0000122E : data <= 8'b00000000 ;
			15'h0000122F : data <= 8'b00000000 ;
			15'h00001230 : data <= 8'b00000000 ;
			15'h00001231 : data <= 8'b00000000 ;
			15'h00001232 : data <= 8'b00000000 ;
			15'h00001233 : data <= 8'b00000000 ;
			15'h00001234 : data <= 8'b00000000 ;
			15'h00001235 : data <= 8'b00000000 ;
			15'h00001236 : data <= 8'b00000000 ;
			15'h00001237 : data <= 8'b00000000 ;
			15'h00001238 : data <= 8'b00000000 ;
			15'h00001239 : data <= 8'b00000000 ;
			15'h0000123A : data <= 8'b00000000 ;
			15'h0000123B : data <= 8'b00000000 ;
			15'h0000123C : data <= 8'b00000000 ;
			15'h0000123D : data <= 8'b00000000 ;
			15'h0000123E : data <= 8'b00000000 ;
			15'h0000123F : data <= 8'b00000000 ;
			15'h00001240 : data <= 8'b00000000 ;
			15'h00001241 : data <= 8'b00000000 ;
			15'h00001242 : data <= 8'b00000000 ;
			15'h00001243 : data <= 8'b00000000 ;
			15'h00001244 : data <= 8'b00000000 ;
			15'h00001245 : data <= 8'b00000000 ;
			15'h00001246 : data <= 8'b00000000 ;
			15'h00001247 : data <= 8'b00000000 ;
			15'h00001248 : data <= 8'b00000000 ;
			15'h00001249 : data <= 8'b00000000 ;
			15'h0000124A : data <= 8'b00000000 ;
			15'h0000124B : data <= 8'b00000000 ;
			15'h0000124C : data <= 8'b00000000 ;
			15'h0000124D : data <= 8'b00000000 ;
			15'h0000124E : data <= 8'b00000000 ;
			15'h0000124F : data <= 8'b00000000 ;
			15'h00001250 : data <= 8'b00000000 ;
			15'h00001251 : data <= 8'b00000000 ;
			15'h00001252 : data <= 8'b00000000 ;
			15'h00001253 : data <= 8'b00000000 ;
			15'h00001254 : data <= 8'b00000000 ;
			15'h00001255 : data <= 8'b00000000 ;
			15'h00001256 : data <= 8'b00000000 ;
			15'h00001257 : data <= 8'b00000000 ;
			15'h00001258 : data <= 8'b00000000 ;
			15'h00001259 : data <= 8'b00000000 ;
			15'h0000125A : data <= 8'b00000000 ;
			15'h0000125B : data <= 8'b00000000 ;
			15'h0000125C : data <= 8'b00000000 ;
			15'h0000125D : data <= 8'b00000000 ;
			15'h0000125E : data <= 8'b00000000 ;
			15'h0000125F : data <= 8'b00000000 ;
			15'h00001260 : data <= 8'b00000000 ;
			15'h00001261 : data <= 8'b00000000 ;
			15'h00001262 : data <= 8'b00000000 ;
			15'h00001263 : data <= 8'b00000000 ;
			15'h00001264 : data <= 8'b00000000 ;
			15'h00001265 : data <= 8'b00000000 ;
			15'h00001266 : data <= 8'b00000000 ;
			15'h00001267 : data <= 8'b00000000 ;
			15'h00001268 : data <= 8'b00000000 ;
			15'h00001269 : data <= 8'b00000000 ;
			15'h0000126A : data <= 8'b00000000 ;
			15'h0000126B : data <= 8'b00000000 ;
			15'h0000126C : data <= 8'b00000000 ;
			15'h0000126D : data <= 8'b00000000 ;
			15'h0000126E : data <= 8'b00000000 ;
			15'h0000126F : data <= 8'b00000000 ;
			15'h00001270 : data <= 8'b00000000 ;
			15'h00001271 : data <= 8'b00000000 ;
			15'h00001272 : data <= 8'b00000000 ;
			15'h00001273 : data <= 8'b00000000 ;
			15'h00001274 : data <= 8'b00000000 ;
			15'h00001275 : data <= 8'b00000000 ;
			15'h00001276 : data <= 8'b00000000 ;
			15'h00001277 : data <= 8'b00000000 ;
			15'h00001278 : data <= 8'b00000000 ;
			15'h00001279 : data <= 8'b00000000 ;
			15'h0000127A : data <= 8'b00000000 ;
			15'h0000127B : data <= 8'b00000000 ;
			15'h0000127C : data <= 8'b00000000 ;
			15'h0000127D : data <= 8'b00000000 ;
			15'h0000127E : data <= 8'b00000000 ;
			15'h0000127F : data <= 8'b00000000 ;
			15'h00001280 : data <= 8'b00000000 ;
			15'h00001281 : data <= 8'b00000000 ;
			15'h00001282 : data <= 8'b00000000 ;
			15'h00001283 : data <= 8'b00000000 ;
			15'h00001284 : data <= 8'b00000000 ;
			15'h00001285 : data <= 8'b00000000 ;
			15'h00001286 : data <= 8'b00000000 ;
			15'h00001287 : data <= 8'b00000000 ;
			15'h00001288 : data <= 8'b00000000 ;
			15'h00001289 : data <= 8'b00000000 ;
			15'h0000128A : data <= 8'b00000000 ;
			15'h0000128B : data <= 8'b00000000 ;
			15'h0000128C : data <= 8'b00000000 ;
			15'h0000128D : data <= 8'b00000000 ;
			15'h0000128E : data <= 8'b00000000 ;
			15'h0000128F : data <= 8'b00000000 ;
			15'h00001290 : data <= 8'b00000000 ;
			15'h00001291 : data <= 8'b00000000 ;
			15'h00001292 : data <= 8'b00000000 ;
			15'h00001293 : data <= 8'b00000000 ;
			15'h00001294 : data <= 8'b00000000 ;
			15'h00001295 : data <= 8'b00000000 ;
			15'h00001296 : data <= 8'b00000000 ;
			15'h00001297 : data <= 8'b00000000 ;
			15'h00001298 : data <= 8'b00000000 ;
			15'h00001299 : data <= 8'b00000000 ;
			15'h0000129A : data <= 8'b00000000 ;
			15'h0000129B : data <= 8'b00000000 ;
			15'h0000129C : data <= 8'b00000000 ;
			15'h0000129D : data <= 8'b00000000 ;
			15'h0000129E : data <= 8'b00000000 ;
			15'h0000129F : data <= 8'b00000000 ;
			15'h000012A0 : data <= 8'b00000000 ;
			15'h000012A1 : data <= 8'b00000000 ;
			15'h000012A2 : data <= 8'b00000000 ;
			15'h000012A3 : data <= 8'b00000000 ;
			15'h000012A4 : data <= 8'b00000000 ;
			15'h000012A5 : data <= 8'b00000000 ;
			15'h000012A6 : data <= 8'b00000000 ;
			15'h000012A7 : data <= 8'b00000000 ;
			15'h000012A8 : data <= 8'b00000000 ;
			15'h000012A9 : data <= 8'b00000000 ;
			15'h000012AA : data <= 8'b00000000 ;
			15'h000012AB : data <= 8'b00000000 ;
			15'h000012AC : data <= 8'b00000000 ;
			15'h000012AD : data <= 8'b00000000 ;
			15'h000012AE : data <= 8'b00000000 ;
			15'h000012AF : data <= 8'b00000000 ;
			15'h000012B0 : data <= 8'b00000000 ;
			15'h000012B1 : data <= 8'b00000000 ;
			15'h000012B2 : data <= 8'b00000000 ;
			15'h000012B3 : data <= 8'b00000000 ;
			15'h000012B4 : data <= 8'b00000000 ;
			15'h000012B5 : data <= 8'b00000000 ;
			15'h000012B6 : data <= 8'b00000000 ;
			15'h000012B7 : data <= 8'b00000000 ;
			15'h000012B8 : data <= 8'b00000000 ;
			15'h000012B9 : data <= 8'b00000000 ;
			15'h000012BA : data <= 8'b00000000 ;
			15'h000012BB : data <= 8'b00000000 ;
			15'h000012BC : data <= 8'b00000000 ;
			15'h000012BD : data <= 8'b00000000 ;
			15'h000012BE : data <= 8'b00000000 ;
			15'h000012BF : data <= 8'b00000000 ;
			15'h000012C0 : data <= 8'b00000000 ;
			15'h000012C1 : data <= 8'b00000000 ;
			15'h000012C2 : data <= 8'b00000000 ;
			15'h000012C3 : data <= 8'b00000000 ;
			15'h000012C4 : data <= 8'b00000000 ;
			15'h000012C5 : data <= 8'b00000000 ;
			15'h000012C6 : data <= 8'b00000000 ;
			15'h000012C7 : data <= 8'b00000000 ;
			15'h000012C8 : data <= 8'b00000000 ;
			15'h000012C9 : data <= 8'b00000000 ;
			15'h000012CA : data <= 8'b00000000 ;
			15'h000012CB : data <= 8'b00000000 ;
			15'h000012CC : data <= 8'b00000000 ;
			15'h000012CD : data <= 8'b00000000 ;
			15'h000012CE : data <= 8'b00000000 ;
			15'h000012CF : data <= 8'b00000000 ;
			15'h000012D0 : data <= 8'b00000000 ;
			15'h000012D1 : data <= 8'b00000000 ;
			15'h000012D2 : data <= 8'b00000000 ;
			15'h000012D3 : data <= 8'b00000000 ;
			15'h000012D4 : data <= 8'b00000000 ;
			15'h000012D5 : data <= 8'b00000000 ;
			15'h000012D6 : data <= 8'b00000000 ;
			15'h000012D7 : data <= 8'b00000000 ;
			15'h000012D8 : data <= 8'b00000000 ;
			15'h000012D9 : data <= 8'b00000000 ;
			15'h000012DA : data <= 8'b00000000 ;
			15'h000012DB : data <= 8'b00000000 ;
			15'h000012DC : data <= 8'b00000000 ;
			15'h000012DD : data <= 8'b00000000 ;
			15'h000012DE : data <= 8'b00000000 ;
			15'h000012DF : data <= 8'b00000000 ;
			15'h000012E0 : data <= 8'b00000000 ;
			15'h000012E1 : data <= 8'b00000000 ;
			15'h000012E2 : data <= 8'b00000000 ;
			15'h000012E3 : data <= 8'b00000000 ;
			15'h000012E4 : data <= 8'b00000000 ;
			15'h000012E5 : data <= 8'b00000000 ;
			15'h000012E6 : data <= 8'b00000000 ;
			15'h000012E7 : data <= 8'b00000000 ;
			15'h000012E8 : data <= 8'b00000000 ;
			15'h000012E9 : data <= 8'b00000000 ;
			15'h000012EA : data <= 8'b00000000 ;
			15'h000012EB : data <= 8'b00000000 ;
			15'h000012EC : data <= 8'b00000000 ;
			15'h000012ED : data <= 8'b00000000 ;
			15'h000012EE : data <= 8'b00000000 ;
			15'h000012EF : data <= 8'b00000000 ;
			15'h000012F0 : data <= 8'b00000000 ;
			15'h000012F1 : data <= 8'b00000000 ;
			15'h000012F2 : data <= 8'b00000000 ;
			15'h000012F3 : data <= 8'b00000000 ;
			15'h000012F4 : data <= 8'b00000000 ;
			15'h000012F5 : data <= 8'b00000000 ;
			15'h000012F6 : data <= 8'b00000000 ;
			15'h000012F7 : data <= 8'b00000000 ;
			15'h000012F8 : data <= 8'b00000000 ;
			15'h000012F9 : data <= 8'b00000000 ;
			15'h000012FA : data <= 8'b00000000 ;
			15'h000012FB : data <= 8'b00000000 ;
			15'h000012FC : data <= 8'b00000000 ;
			15'h000012FD : data <= 8'b00000000 ;
			15'h000012FE : data <= 8'b00000000 ;
			15'h000012FF : data <= 8'b00000000 ;
			15'h00001300 : data <= 8'b00000000 ;
			15'h00001301 : data <= 8'b00000000 ;
			15'h00001302 : data <= 8'b00000000 ;
			15'h00001303 : data <= 8'b00000000 ;
			15'h00001304 : data <= 8'b00000000 ;
			15'h00001305 : data <= 8'b00000000 ;
			15'h00001306 : data <= 8'b00000000 ;
			15'h00001307 : data <= 8'b00000000 ;
			15'h00001308 : data <= 8'b00000000 ;
			15'h00001309 : data <= 8'b00000000 ;
			15'h0000130A : data <= 8'b00000000 ;
			15'h0000130B : data <= 8'b00000000 ;
			15'h0000130C : data <= 8'b00000000 ;
			15'h0000130D : data <= 8'b00000000 ;
			15'h0000130E : data <= 8'b00000000 ;
			15'h0000130F : data <= 8'b00000000 ;
			15'h00001310 : data <= 8'b00000000 ;
			15'h00001311 : data <= 8'b00000000 ;
			15'h00001312 : data <= 8'b00000000 ;
			15'h00001313 : data <= 8'b00000000 ;
			15'h00001314 : data <= 8'b00000000 ;
			15'h00001315 : data <= 8'b00000000 ;
			15'h00001316 : data <= 8'b00000000 ;
			15'h00001317 : data <= 8'b00000000 ;
			15'h00001318 : data <= 8'b00000000 ;
			15'h00001319 : data <= 8'b00000000 ;
			15'h0000131A : data <= 8'b00000000 ;
			15'h0000131B : data <= 8'b00000000 ;
			15'h0000131C : data <= 8'b00000000 ;
			15'h0000131D : data <= 8'b00000000 ;
			15'h0000131E : data <= 8'b00000000 ;
			15'h0000131F : data <= 8'b00000000 ;
			15'h00001320 : data <= 8'b00000000 ;
			15'h00001321 : data <= 8'b00000000 ;
			15'h00001322 : data <= 8'b00000000 ;
			15'h00001323 : data <= 8'b00000000 ;
			15'h00001324 : data <= 8'b00000000 ;
			15'h00001325 : data <= 8'b00000000 ;
			15'h00001326 : data <= 8'b00000000 ;
			15'h00001327 : data <= 8'b00000000 ;
			15'h00001328 : data <= 8'b00000000 ;
			15'h00001329 : data <= 8'b00000000 ;
			15'h0000132A : data <= 8'b00000000 ;
			15'h0000132B : data <= 8'b00000000 ;
			15'h0000132C : data <= 8'b00000000 ;
			15'h0000132D : data <= 8'b00000000 ;
			15'h0000132E : data <= 8'b00000000 ;
			15'h0000132F : data <= 8'b00000000 ;
			15'h00001330 : data <= 8'b00000000 ;
			15'h00001331 : data <= 8'b00000000 ;
			15'h00001332 : data <= 8'b00000000 ;
			15'h00001333 : data <= 8'b00000000 ;
			15'h00001334 : data <= 8'b00000000 ;
			15'h00001335 : data <= 8'b00000000 ;
			15'h00001336 : data <= 8'b00000000 ;
			15'h00001337 : data <= 8'b00000000 ;
			15'h00001338 : data <= 8'b00000000 ;
			15'h00001339 : data <= 8'b00000000 ;
			15'h0000133A : data <= 8'b00000000 ;
			15'h0000133B : data <= 8'b00000000 ;
			15'h0000133C : data <= 8'b00000000 ;
			15'h0000133D : data <= 8'b00000000 ;
			15'h0000133E : data <= 8'b00000000 ;
			15'h0000133F : data <= 8'b00000000 ;
			15'h00001340 : data <= 8'b00000000 ;
			15'h00001341 : data <= 8'b00000000 ;
			15'h00001342 : data <= 8'b00000000 ;
			15'h00001343 : data <= 8'b00000000 ;
			15'h00001344 : data <= 8'b00000000 ;
			15'h00001345 : data <= 8'b00000000 ;
			15'h00001346 : data <= 8'b00000000 ;
			15'h00001347 : data <= 8'b00000000 ;
			15'h00001348 : data <= 8'b00000000 ;
			15'h00001349 : data <= 8'b00000000 ;
			15'h0000134A : data <= 8'b00000000 ;
			15'h0000134B : data <= 8'b00000000 ;
			15'h0000134C : data <= 8'b00000000 ;
			15'h0000134D : data <= 8'b00000000 ;
			15'h0000134E : data <= 8'b00000000 ;
			15'h0000134F : data <= 8'b00000000 ;
			15'h00001350 : data <= 8'b00000000 ;
			15'h00001351 : data <= 8'b00000000 ;
			15'h00001352 : data <= 8'b00000000 ;
			15'h00001353 : data <= 8'b00000000 ;
			15'h00001354 : data <= 8'b00000000 ;
			15'h00001355 : data <= 8'b00000000 ;
			15'h00001356 : data <= 8'b00000000 ;
			15'h00001357 : data <= 8'b00000000 ;
			15'h00001358 : data <= 8'b00000000 ;
			15'h00001359 : data <= 8'b00000000 ;
			15'h0000135A : data <= 8'b00000000 ;
			15'h0000135B : data <= 8'b00000000 ;
			15'h0000135C : data <= 8'b00000000 ;
			15'h0000135D : data <= 8'b00000000 ;
			15'h0000135E : data <= 8'b00000000 ;
			15'h0000135F : data <= 8'b00000000 ;
			15'h00001360 : data <= 8'b00000000 ;
			15'h00001361 : data <= 8'b00000000 ;
			15'h00001362 : data <= 8'b00000000 ;
			15'h00001363 : data <= 8'b00000000 ;
			15'h00001364 : data <= 8'b00000000 ;
			15'h00001365 : data <= 8'b00000000 ;
			15'h00001366 : data <= 8'b00000000 ;
			15'h00001367 : data <= 8'b00000000 ;
			15'h00001368 : data <= 8'b00000000 ;
			15'h00001369 : data <= 8'b00000000 ;
			15'h0000136A : data <= 8'b00000000 ;
			15'h0000136B : data <= 8'b00000000 ;
			15'h0000136C : data <= 8'b00000000 ;
			15'h0000136D : data <= 8'b00000000 ;
			15'h0000136E : data <= 8'b00000000 ;
			15'h0000136F : data <= 8'b00000000 ;
			15'h00001370 : data <= 8'b00000000 ;
			15'h00001371 : data <= 8'b00000000 ;
			15'h00001372 : data <= 8'b00000000 ;
			15'h00001373 : data <= 8'b00000000 ;
			15'h00001374 : data <= 8'b00000000 ;
			15'h00001375 : data <= 8'b00000000 ;
			15'h00001376 : data <= 8'b00000000 ;
			15'h00001377 : data <= 8'b00000000 ;
			15'h00001378 : data <= 8'b00000000 ;
			15'h00001379 : data <= 8'b00000000 ;
			15'h0000137A : data <= 8'b00000000 ;
			15'h0000137B : data <= 8'b00000000 ;
			15'h0000137C : data <= 8'b00000000 ;
			15'h0000137D : data <= 8'b00000000 ;
			15'h0000137E : data <= 8'b00000000 ;
			15'h0000137F : data <= 8'b00000000 ;
			15'h00001380 : data <= 8'b00000000 ;
			15'h00001381 : data <= 8'b00000000 ;
			15'h00001382 : data <= 8'b00000000 ;
			15'h00001383 : data <= 8'b00000000 ;
			15'h00001384 : data <= 8'b00000000 ;
			15'h00001385 : data <= 8'b00000000 ;
			15'h00001386 : data <= 8'b00000000 ;
			15'h00001387 : data <= 8'b00000000 ;
			15'h00001388 : data <= 8'b00000000 ;
			15'h00001389 : data <= 8'b00000000 ;
			15'h0000138A : data <= 8'b00000000 ;
			15'h0000138B : data <= 8'b00000000 ;
			15'h0000138C : data <= 8'b00000000 ;
			15'h0000138D : data <= 8'b00000000 ;
			15'h0000138E : data <= 8'b00000000 ;
			15'h0000138F : data <= 8'b00000000 ;
			15'h00001390 : data <= 8'b00000000 ;
			15'h00001391 : data <= 8'b00000000 ;
			15'h00001392 : data <= 8'b00000000 ;
			15'h00001393 : data <= 8'b00000000 ;
			15'h00001394 : data <= 8'b00000000 ;
			15'h00001395 : data <= 8'b00000000 ;
			15'h00001396 : data <= 8'b00000000 ;
			15'h00001397 : data <= 8'b00000000 ;
			15'h00001398 : data <= 8'b00000000 ;
			15'h00001399 : data <= 8'b00000000 ;
			15'h0000139A : data <= 8'b00000000 ;
			15'h0000139B : data <= 8'b00000000 ;
			15'h0000139C : data <= 8'b00000000 ;
			15'h0000139D : data <= 8'b00000000 ;
			15'h0000139E : data <= 8'b00000000 ;
			15'h0000139F : data <= 8'b00000000 ;
			15'h000013A0 : data <= 8'b00000000 ;
			15'h000013A1 : data <= 8'b00000000 ;
			15'h000013A2 : data <= 8'b00000000 ;
			15'h000013A3 : data <= 8'b00000000 ;
			15'h000013A4 : data <= 8'b00000000 ;
			15'h000013A5 : data <= 8'b00000000 ;
			15'h000013A6 : data <= 8'b00000000 ;
			15'h000013A7 : data <= 8'b00000000 ;
			15'h000013A8 : data <= 8'b00000000 ;
			15'h000013A9 : data <= 8'b00000000 ;
			15'h000013AA : data <= 8'b00000000 ;
			15'h000013AB : data <= 8'b00000000 ;
			15'h000013AC : data <= 8'b00000000 ;
			15'h000013AD : data <= 8'b00000000 ;
			15'h000013AE : data <= 8'b00000000 ;
			15'h000013AF : data <= 8'b00000000 ;
			15'h000013B0 : data <= 8'b00000000 ;
			15'h000013B1 : data <= 8'b00000000 ;
			15'h000013B2 : data <= 8'b00000000 ;
			15'h000013B3 : data <= 8'b00000000 ;
			15'h000013B4 : data <= 8'b00000000 ;
			15'h000013B5 : data <= 8'b00000000 ;
			15'h000013B6 : data <= 8'b00000000 ;
			15'h000013B7 : data <= 8'b00000000 ;
			15'h000013B8 : data <= 8'b00000000 ;
			15'h000013B9 : data <= 8'b00000000 ;
			15'h000013BA : data <= 8'b00000000 ;
			15'h000013BB : data <= 8'b00000000 ;
			15'h000013BC : data <= 8'b00000000 ;
			15'h000013BD : data <= 8'b00000000 ;
			15'h000013BE : data <= 8'b00000000 ;
			15'h000013BF : data <= 8'b00000000 ;
			15'h000013C0 : data <= 8'b00000000 ;
			15'h000013C1 : data <= 8'b00000000 ;
			15'h000013C2 : data <= 8'b00000000 ;
			15'h000013C3 : data <= 8'b00000000 ;
			15'h000013C4 : data <= 8'b00000000 ;
			15'h000013C5 : data <= 8'b00000000 ;
			15'h000013C6 : data <= 8'b00000000 ;
			15'h000013C7 : data <= 8'b00000000 ;
			15'h000013C8 : data <= 8'b00000000 ;
			15'h000013C9 : data <= 8'b00000000 ;
			15'h000013CA : data <= 8'b00000000 ;
			15'h000013CB : data <= 8'b00000000 ;
			15'h000013CC : data <= 8'b00000000 ;
			15'h000013CD : data <= 8'b00000000 ;
			15'h000013CE : data <= 8'b00000000 ;
			15'h000013CF : data <= 8'b00000000 ;
			15'h000013D0 : data <= 8'b00000000 ;
			15'h000013D1 : data <= 8'b00000000 ;
			15'h000013D2 : data <= 8'b00000000 ;
			15'h000013D3 : data <= 8'b00000000 ;
			15'h000013D4 : data <= 8'b00000000 ;
			15'h000013D5 : data <= 8'b00000000 ;
			15'h000013D6 : data <= 8'b00000000 ;
			15'h000013D7 : data <= 8'b00000000 ;
			15'h000013D8 : data <= 8'b00000000 ;
			15'h000013D9 : data <= 8'b00000000 ;
			15'h000013DA : data <= 8'b00000000 ;
			15'h000013DB : data <= 8'b00000000 ;
			15'h000013DC : data <= 8'b00000000 ;
			15'h000013DD : data <= 8'b00000000 ;
			15'h000013DE : data <= 8'b00000000 ;
			15'h000013DF : data <= 8'b00000000 ;
			15'h000013E0 : data <= 8'b00000000 ;
			15'h000013E1 : data <= 8'b00000000 ;
			15'h000013E2 : data <= 8'b00000000 ;
			15'h000013E3 : data <= 8'b00000000 ;
			15'h000013E4 : data <= 8'b00000000 ;
			15'h000013E5 : data <= 8'b00000000 ;
			15'h000013E6 : data <= 8'b00000000 ;
			15'h000013E7 : data <= 8'b00000000 ;
			15'h000013E8 : data <= 8'b00000000 ;
			15'h000013E9 : data <= 8'b00000000 ;
			15'h000013EA : data <= 8'b00000000 ;
			15'h000013EB : data <= 8'b00000000 ;
			15'h000013EC : data <= 8'b00000000 ;
			15'h000013ED : data <= 8'b00000000 ;
			15'h000013EE : data <= 8'b00000000 ;
			15'h000013EF : data <= 8'b00000000 ;
			15'h000013F0 : data <= 8'b00000000 ;
			15'h000013F1 : data <= 8'b00000000 ;
			15'h000013F2 : data <= 8'b00000000 ;
			15'h000013F3 : data <= 8'b00000000 ;
			15'h000013F4 : data <= 8'b00000000 ;
			15'h000013F5 : data <= 8'b00000000 ;
			15'h000013F6 : data <= 8'b00000000 ;
			15'h000013F7 : data <= 8'b00000000 ;
			15'h000013F8 : data <= 8'b00000000 ;
			15'h000013F9 : data <= 8'b00000000 ;
			15'h000013FA : data <= 8'b00000000 ;
			15'h000013FB : data <= 8'b00000000 ;
			15'h000013FC : data <= 8'b00000000 ;
			15'h000013FD : data <= 8'b00000000 ;
			15'h000013FE : data <= 8'b00000000 ;
			15'h000013FF : data <= 8'b00000000 ;
			15'h00001400 : data <= 8'b00000000 ;
			15'h00001401 : data <= 8'b00000000 ;
			15'h00001402 : data <= 8'b00000000 ;
			15'h00001403 : data <= 8'b00000000 ;
			15'h00001404 : data <= 8'b00000000 ;
			15'h00001405 : data <= 8'b00000000 ;
			15'h00001406 : data <= 8'b00000000 ;
			15'h00001407 : data <= 8'b00000000 ;
			15'h00001408 : data <= 8'b00000000 ;
			15'h00001409 : data <= 8'b00000000 ;
			15'h0000140A : data <= 8'b00000000 ;
			15'h0000140B : data <= 8'b00000000 ;
			15'h0000140C : data <= 8'b00000000 ;
			15'h0000140D : data <= 8'b00000000 ;
			15'h0000140E : data <= 8'b00000000 ;
			15'h0000140F : data <= 8'b00000000 ;
			15'h00001410 : data <= 8'b00000000 ;
			15'h00001411 : data <= 8'b00000000 ;
			15'h00001412 : data <= 8'b00000000 ;
			15'h00001413 : data <= 8'b00000000 ;
			15'h00001414 : data <= 8'b00000000 ;
			15'h00001415 : data <= 8'b00000000 ;
			15'h00001416 : data <= 8'b00000000 ;
			15'h00001417 : data <= 8'b00000000 ;
			15'h00001418 : data <= 8'b00000000 ;
			15'h00001419 : data <= 8'b00000000 ;
			15'h0000141A : data <= 8'b00000000 ;
			15'h0000141B : data <= 8'b00000000 ;
			15'h0000141C : data <= 8'b00000000 ;
			15'h0000141D : data <= 8'b00000000 ;
			15'h0000141E : data <= 8'b00000000 ;
			15'h0000141F : data <= 8'b00000000 ;
			15'h00001420 : data <= 8'b00000000 ;
			15'h00001421 : data <= 8'b00000000 ;
			15'h00001422 : data <= 8'b00000000 ;
			15'h00001423 : data <= 8'b00000000 ;
			15'h00001424 : data <= 8'b00000000 ;
			15'h00001425 : data <= 8'b00000000 ;
			15'h00001426 : data <= 8'b00000000 ;
			15'h00001427 : data <= 8'b00000000 ;
			15'h00001428 : data <= 8'b00000000 ;
			15'h00001429 : data <= 8'b00000000 ;
			15'h0000142A : data <= 8'b00000000 ;
			15'h0000142B : data <= 8'b00000000 ;
			15'h0000142C : data <= 8'b00000000 ;
			15'h0000142D : data <= 8'b00000000 ;
			15'h0000142E : data <= 8'b00000000 ;
			15'h0000142F : data <= 8'b00000000 ;
			15'h00001430 : data <= 8'b00000000 ;
			15'h00001431 : data <= 8'b00000000 ;
			15'h00001432 : data <= 8'b00000000 ;
			15'h00001433 : data <= 8'b00000000 ;
			15'h00001434 : data <= 8'b00000000 ;
			15'h00001435 : data <= 8'b00000000 ;
			15'h00001436 : data <= 8'b00000000 ;
			15'h00001437 : data <= 8'b00000000 ;
			15'h00001438 : data <= 8'b00000000 ;
			15'h00001439 : data <= 8'b00000000 ;
			15'h0000143A : data <= 8'b00000000 ;
			15'h0000143B : data <= 8'b00000000 ;
			15'h0000143C : data <= 8'b00000000 ;
			15'h0000143D : data <= 8'b00000000 ;
			15'h0000143E : data <= 8'b00000000 ;
			15'h0000143F : data <= 8'b00000000 ;
			15'h00001440 : data <= 8'b00000000 ;
			15'h00001441 : data <= 8'b00000000 ;
			15'h00001442 : data <= 8'b00000000 ;
			15'h00001443 : data <= 8'b00000000 ;
			15'h00001444 : data <= 8'b00000000 ;
			15'h00001445 : data <= 8'b00000000 ;
			15'h00001446 : data <= 8'b00000000 ;
			15'h00001447 : data <= 8'b00000000 ;
			15'h00001448 : data <= 8'b00000000 ;
			15'h00001449 : data <= 8'b00000000 ;
			15'h0000144A : data <= 8'b00000000 ;
			15'h0000144B : data <= 8'b00000000 ;
			15'h0000144C : data <= 8'b00000000 ;
			15'h0000144D : data <= 8'b00000000 ;
			15'h0000144E : data <= 8'b00000000 ;
			15'h0000144F : data <= 8'b00000000 ;
			15'h00001450 : data <= 8'b00000000 ;
			15'h00001451 : data <= 8'b00000000 ;
			15'h00001452 : data <= 8'b00000000 ;
			15'h00001453 : data <= 8'b00000000 ;
			15'h00001454 : data <= 8'b00000000 ;
			15'h00001455 : data <= 8'b00000000 ;
			15'h00001456 : data <= 8'b00000000 ;
			15'h00001457 : data <= 8'b00000000 ;
			15'h00001458 : data <= 8'b00000000 ;
			15'h00001459 : data <= 8'b00000000 ;
			15'h0000145A : data <= 8'b00000000 ;
			15'h0000145B : data <= 8'b00000000 ;
			15'h0000145C : data <= 8'b00000000 ;
			15'h0000145D : data <= 8'b00000000 ;
			15'h0000145E : data <= 8'b00000000 ;
			15'h0000145F : data <= 8'b00000000 ;
			15'h00001460 : data <= 8'b00000000 ;
			15'h00001461 : data <= 8'b00000000 ;
			15'h00001462 : data <= 8'b00000000 ;
			15'h00001463 : data <= 8'b00000000 ;
			15'h00001464 : data <= 8'b00000000 ;
			15'h00001465 : data <= 8'b00000000 ;
			15'h00001466 : data <= 8'b00000000 ;
			15'h00001467 : data <= 8'b00000000 ;
			15'h00001468 : data <= 8'b00000000 ;
			15'h00001469 : data <= 8'b00000000 ;
			15'h0000146A : data <= 8'b00000000 ;
			15'h0000146B : data <= 8'b00000000 ;
			15'h0000146C : data <= 8'b00000000 ;
			15'h0000146D : data <= 8'b00000000 ;
			15'h0000146E : data <= 8'b00000000 ;
			15'h0000146F : data <= 8'b00000000 ;
			15'h00001470 : data <= 8'b00000000 ;
			15'h00001471 : data <= 8'b00000000 ;
			15'h00001472 : data <= 8'b00000000 ;
			15'h00001473 : data <= 8'b00000000 ;
			15'h00001474 : data <= 8'b00000000 ;
			15'h00001475 : data <= 8'b00000000 ;
			15'h00001476 : data <= 8'b00000000 ;
			15'h00001477 : data <= 8'b00000000 ;
			15'h00001478 : data <= 8'b00000000 ;
			15'h00001479 : data <= 8'b00000000 ;
			15'h0000147A : data <= 8'b00000000 ;
			15'h0000147B : data <= 8'b00000000 ;
			15'h0000147C : data <= 8'b00000000 ;
			15'h0000147D : data <= 8'b00000000 ;
			15'h0000147E : data <= 8'b00000000 ;
			15'h0000147F : data <= 8'b00000000 ;
			15'h00001480 : data <= 8'b00000000 ;
			15'h00001481 : data <= 8'b00000000 ;
			15'h00001482 : data <= 8'b00000000 ;
			15'h00001483 : data <= 8'b00000000 ;
			15'h00001484 : data <= 8'b00000000 ;
			15'h00001485 : data <= 8'b00000000 ;
			15'h00001486 : data <= 8'b00000000 ;
			15'h00001487 : data <= 8'b00000000 ;
			15'h00001488 : data <= 8'b00000000 ;
			15'h00001489 : data <= 8'b00000000 ;
			15'h0000148A : data <= 8'b00000000 ;
			15'h0000148B : data <= 8'b00000000 ;
			15'h0000148C : data <= 8'b00000000 ;
			15'h0000148D : data <= 8'b00000000 ;
			15'h0000148E : data <= 8'b00000000 ;
			15'h0000148F : data <= 8'b00000000 ;
			15'h00001490 : data <= 8'b00000000 ;
			15'h00001491 : data <= 8'b00000000 ;
			15'h00001492 : data <= 8'b00000000 ;
			15'h00001493 : data <= 8'b00000000 ;
			15'h00001494 : data <= 8'b00000000 ;
			15'h00001495 : data <= 8'b00000000 ;
			15'h00001496 : data <= 8'b00000000 ;
			15'h00001497 : data <= 8'b00000000 ;
			15'h00001498 : data <= 8'b00000000 ;
			15'h00001499 : data <= 8'b00000000 ;
			15'h0000149A : data <= 8'b00000000 ;
			15'h0000149B : data <= 8'b00000000 ;
			15'h0000149C : data <= 8'b00000000 ;
			15'h0000149D : data <= 8'b00000000 ;
			15'h0000149E : data <= 8'b00000000 ;
			15'h0000149F : data <= 8'b00000000 ;
			15'h000014A0 : data <= 8'b00000000 ;
			15'h000014A1 : data <= 8'b00000000 ;
			15'h000014A2 : data <= 8'b00000000 ;
			15'h000014A3 : data <= 8'b00000000 ;
			15'h000014A4 : data <= 8'b00000000 ;
			15'h000014A5 : data <= 8'b00000000 ;
			15'h000014A6 : data <= 8'b00000000 ;
			15'h000014A7 : data <= 8'b00000000 ;
			15'h000014A8 : data <= 8'b00000000 ;
			15'h000014A9 : data <= 8'b00000000 ;
			15'h000014AA : data <= 8'b00000000 ;
			15'h000014AB : data <= 8'b00000000 ;
			15'h000014AC : data <= 8'b00000000 ;
			15'h000014AD : data <= 8'b00000000 ;
			15'h000014AE : data <= 8'b00000000 ;
			15'h000014AF : data <= 8'b00000000 ;
			15'h000014B0 : data <= 8'b00000000 ;
			15'h000014B1 : data <= 8'b00000000 ;
			15'h000014B2 : data <= 8'b00000000 ;
			15'h000014B3 : data <= 8'b00000000 ;
			15'h000014B4 : data <= 8'b00000000 ;
			15'h000014B5 : data <= 8'b00000000 ;
			15'h000014B6 : data <= 8'b00000000 ;
			15'h000014B7 : data <= 8'b00000000 ;
			15'h000014B8 : data <= 8'b00000000 ;
			15'h000014B9 : data <= 8'b00000000 ;
			15'h000014BA : data <= 8'b00000000 ;
			15'h000014BB : data <= 8'b00000000 ;
			15'h000014BC : data <= 8'b00000000 ;
			15'h000014BD : data <= 8'b00000000 ;
			15'h000014BE : data <= 8'b00000000 ;
			15'h000014BF : data <= 8'b00000000 ;
			15'h000014C0 : data <= 8'b00000000 ;
			15'h000014C1 : data <= 8'b00000000 ;
			15'h000014C2 : data <= 8'b00000000 ;
			15'h000014C3 : data <= 8'b00000000 ;
			15'h000014C4 : data <= 8'b00000000 ;
			15'h000014C5 : data <= 8'b00000000 ;
			15'h000014C6 : data <= 8'b00000000 ;
			15'h000014C7 : data <= 8'b00000000 ;
			15'h000014C8 : data <= 8'b00000000 ;
			15'h000014C9 : data <= 8'b00000000 ;
			15'h000014CA : data <= 8'b00000000 ;
			15'h000014CB : data <= 8'b00000000 ;
			15'h000014CC : data <= 8'b00000000 ;
			15'h000014CD : data <= 8'b00000000 ;
			15'h000014CE : data <= 8'b00000000 ;
			15'h000014CF : data <= 8'b00000000 ;
			15'h000014D0 : data <= 8'b00000000 ;
			15'h000014D1 : data <= 8'b00000000 ;
			15'h000014D2 : data <= 8'b00000000 ;
			15'h000014D3 : data <= 8'b00000000 ;
			15'h000014D4 : data <= 8'b00000000 ;
			15'h000014D5 : data <= 8'b00000000 ;
			15'h000014D6 : data <= 8'b00000000 ;
			15'h000014D7 : data <= 8'b00000000 ;
			15'h000014D8 : data <= 8'b00000000 ;
			15'h000014D9 : data <= 8'b00000000 ;
			15'h000014DA : data <= 8'b00000000 ;
			15'h000014DB : data <= 8'b00000000 ;
			15'h000014DC : data <= 8'b00000000 ;
			15'h000014DD : data <= 8'b00000000 ;
			15'h000014DE : data <= 8'b00000000 ;
			15'h000014DF : data <= 8'b00000000 ;
			15'h000014E0 : data <= 8'b00000000 ;
			15'h000014E1 : data <= 8'b00000000 ;
			15'h000014E2 : data <= 8'b00000000 ;
			15'h000014E3 : data <= 8'b00000000 ;
			15'h000014E4 : data <= 8'b00000000 ;
			15'h000014E5 : data <= 8'b00000000 ;
			15'h000014E6 : data <= 8'b00000000 ;
			15'h000014E7 : data <= 8'b00000000 ;
			15'h000014E8 : data <= 8'b00000000 ;
			15'h000014E9 : data <= 8'b00000000 ;
			15'h000014EA : data <= 8'b00000000 ;
			15'h000014EB : data <= 8'b00000000 ;
			15'h000014EC : data <= 8'b00000000 ;
			15'h000014ED : data <= 8'b00000000 ;
			15'h000014EE : data <= 8'b00000000 ;
			15'h000014EF : data <= 8'b00000000 ;
			15'h000014F0 : data <= 8'b00000000 ;
			15'h000014F1 : data <= 8'b00000000 ;
			15'h000014F2 : data <= 8'b00000000 ;
			15'h000014F3 : data <= 8'b00000000 ;
			15'h000014F4 : data <= 8'b00000000 ;
			15'h000014F5 : data <= 8'b00000000 ;
			15'h000014F6 : data <= 8'b00000000 ;
			15'h000014F7 : data <= 8'b00000000 ;
			15'h000014F8 : data <= 8'b00000000 ;
			15'h000014F9 : data <= 8'b00000000 ;
			15'h000014FA : data <= 8'b00000000 ;
			15'h000014FB : data <= 8'b00000000 ;
			15'h000014FC : data <= 8'b00000000 ;
			15'h000014FD : data <= 8'b00000000 ;
			15'h000014FE : data <= 8'b00000000 ;
			15'h000014FF : data <= 8'b00000000 ;
			15'h00001500 : data <= 8'b00000000 ;
			15'h00001501 : data <= 8'b00000000 ;
			15'h00001502 : data <= 8'b00000000 ;
			15'h00001503 : data <= 8'b00000000 ;
			15'h00001504 : data <= 8'b00000000 ;
			15'h00001505 : data <= 8'b00000000 ;
			15'h00001506 : data <= 8'b00000000 ;
			15'h00001507 : data <= 8'b00000000 ;
			15'h00001508 : data <= 8'b00000000 ;
			15'h00001509 : data <= 8'b00000000 ;
			15'h0000150A : data <= 8'b00000000 ;
			15'h0000150B : data <= 8'b00000000 ;
			15'h0000150C : data <= 8'b00000000 ;
			15'h0000150D : data <= 8'b00000000 ;
			15'h0000150E : data <= 8'b00000000 ;
			15'h0000150F : data <= 8'b00000000 ;
			15'h00001510 : data <= 8'b00000000 ;
			15'h00001511 : data <= 8'b00000000 ;
			15'h00001512 : data <= 8'b00000000 ;
			15'h00001513 : data <= 8'b00000000 ;
			15'h00001514 : data <= 8'b00000000 ;
			15'h00001515 : data <= 8'b00000000 ;
			15'h00001516 : data <= 8'b00000000 ;
			15'h00001517 : data <= 8'b00000000 ;
			15'h00001518 : data <= 8'b00000000 ;
			15'h00001519 : data <= 8'b00000000 ;
			15'h0000151A : data <= 8'b00000000 ;
			15'h0000151B : data <= 8'b00000000 ;
			15'h0000151C : data <= 8'b00000000 ;
			15'h0000151D : data <= 8'b00000000 ;
			15'h0000151E : data <= 8'b00000000 ;
			15'h0000151F : data <= 8'b00000000 ;
			15'h00001520 : data <= 8'b00000000 ;
			15'h00001521 : data <= 8'b00000000 ;
			15'h00001522 : data <= 8'b00000000 ;
			15'h00001523 : data <= 8'b00000000 ;
			15'h00001524 : data <= 8'b00000000 ;
			15'h00001525 : data <= 8'b00000000 ;
			15'h00001526 : data <= 8'b00000000 ;
			15'h00001527 : data <= 8'b00000000 ;
			15'h00001528 : data <= 8'b00000000 ;
			15'h00001529 : data <= 8'b00000000 ;
			15'h0000152A : data <= 8'b00000000 ;
			15'h0000152B : data <= 8'b00000000 ;
			15'h0000152C : data <= 8'b00000000 ;
			15'h0000152D : data <= 8'b00000000 ;
			15'h0000152E : data <= 8'b00000000 ;
			15'h0000152F : data <= 8'b00000000 ;
			15'h00001530 : data <= 8'b00000000 ;
			15'h00001531 : data <= 8'b00000000 ;
			15'h00001532 : data <= 8'b00000000 ;
			15'h00001533 : data <= 8'b00000000 ;
			15'h00001534 : data <= 8'b00000000 ;
			15'h00001535 : data <= 8'b00000000 ;
			15'h00001536 : data <= 8'b00000000 ;
			15'h00001537 : data <= 8'b00000000 ;
			15'h00001538 : data <= 8'b00000000 ;
			15'h00001539 : data <= 8'b00000000 ;
			15'h0000153A : data <= 8'b00000000 ;
			15'h0000153B : data <= 8'b00000000 ;
			15'h0000153C : data <= 8'b00000000 ;
			15'h0000153D : data <= 8'b00000000 ;
			15'h0000153E : data <= 8'b00000000 ;
			15'h0000153F : data <= 8'b00000000 ;
			15'h00001540 : data <= 8'b00000000 ;
			15'h00001541 : data <= 8'b00000000 ;
			15'h00001542 : data <= 8'b00000000 ;
			15'h00001543 : data <= 8'b00000000 ;
			15'h00001544 : data <= 8'b00000000 ;
			15'h00001545 : data <= 8'b00000000 ;
			15'h00001546 : data <= 8'b00000000 ;
			15'h00001547 : data <= 8'b00000000 ;
			15'h00001548 : data <= 8'b00000000 ;
			15'h00001549 : data <= 8'b00000000 ;
			15'h0000154A : data <= 8'b00000000 ;
			15'h0000154B : data <= 8'b00000000 ;
			15'h0000154C : data <= 8'b00000000 ;
			15'h0000154D : data <= 8'b00000000 ;
			15'h0000154E : data <= 8'b00000000 ;
			15'h0000154F : data <= 8'b00000000 ;
			15'h00001550 : data <= 8'b00000000 ;
			15'h00001551 : data <= 8'b00000000 ;
			15'h00001552 : data <= 8'b00000000 ;
			15'h00001553 : data <= 8'b00000000 ;
			15'h00001554 : data <= 8'b00000000 ;
			15'h00001555 : data <= 8'b00000000 ;
			15'h00001556 : data <= 8'b00000000 ;
			15'h00001557 : data <= 8'b00000000 ;
			15'h00001558 : data <= 8'b00000000 ;
			15'h00001559 : data <= 8'b00000000 ;
			15'h0000155A : data <= 8'b00000000 ;
			15'h0000155B : data <= 8'b00000000 ;
			15'h0000155C : data <= 8'b00000000 ;
			15'h0000155D : data <= 8'b00000000 ;
			15'h0000155E : data <= 8'b00000000 ;
			15'h0000155F : data <= 8'b00000000 ;
			15'h00001560 : data <= 8'b00000000 ;
			15'h00001561 : data <= 8'b00000000 ;
			15'h00001562 : data <= 8'b00000000 ;
			15'h00001563 : data <= 8'b00000000 ;
			15'h00001564 : data <= 8'b00000000 ;
			15'h00001565 : data <= 8'b00000000 ;
			15'h00001566 : data <= 8'b00000000 ;
			15'h00001567 : data <= 8'b00000000 ;
			15'h00001568 : data <= 8'b00000000 ;
			15'h00001569 : data <= 8'b00000000 ;
			15'h0000156A : data <= 8'b00000000 ;
			15'h0000156B : data <= 8'b00000000 ;
			15'h0000156C : data <= 8'b00000000 ;
			15'h0000156D : data <= 8'b00000000 ;
			15'h0000156E : data <= 8'b00000000 ;
			15'h0000156F : data <= 8'b00000000 ;
			15'h00001570 : data <= 8'b00000000 ;
			15'h00001571 : data <= 8'b00000000 ;
			15'h00001572 : data <= 8'b00000000 ;
			15'h00001573 : data <= 8'b00000000 ;
			15'h00001574 : data <= 8'b00000000 ;
			15'h00001575 : data <= 8'b00000000 ;
			15'h00001576 : data <= 8'b00000000 ;
			15'h00001577 : data <= 8'b00000000 ;
			15'h00001578 : data <= 8'b00000000 ;
			15'h00001579 : data <= 8'b00000000 ;
			15'h0000157A : data <= 8'b00000000 ;
			15'h0000157B : data <= 8'b00000000 ;
			15'h0000157C : data <= 8'b00000000 ;
			15'h0000157D : data <= 8'b00000000 ;
			15'h0000157E : data <= 8'b00000000 ;
			15'h0000157F : data <= 8'b00000000 ;
			15'h00001580 : data <= 8'b00000000 ;
			15'h00001581 : data <= 8'b00000000 ;
			15'h00001582 : data <= 8'b00000000 ;
			15'h00001583 : data <= 8'b00000000 ;
			15'h00001584 : data <= 8'b00000000 ;
			15'h00001585 : data <= 8'b00000000 ;
			15'h00001586 : data <= 8'b00000000 ;
			15'h00001587 : data <= 8'b00000000 ;
			15'h00001588 : data <= 8'b00000000 ;
			15'h00001589 : data <= 8'b00000000 ;
			15'h0000158A : data <= 8'b00000000 ;
			15'h0000158B : data <= 8'b00000000 ;
			15'h0000158C : data <= 8'b00000000 ;
			15'h0000158D : data <= 8'b00000000 ;
			15'h0000158E : data <= 8'b00000000 ;
			15'h0000158F : data <= 8'b00000000 ;
			15'h00001590 : data <= 8'b00000000 ;
			15'h00001591 : data <= 8'b00000000 ;
			15'h00001592 : data <= 8'b00000000 ;
			15'h00001593 : data <= 8'b00000000 ;
			15'h00001594 : data <= 8'b00000000 ;
			15'h00001595 : data <= 8'b00000000 ;
			15'h00001596 : data <= 8'b00000000 ;
			15'h00001597 : data <= 8'b00000000 ;
			15'h00001598 : data <= 8'b00000000 ;
			15'h00001599 : data <= 8'b00000000 ;
			15'h0000159A : data <= 8'b00000000 ;
			15'h0000159B : data <= 8'b00000000 ;
			15'h0000159C : data <= 8'b00000000 ;
			15'h0000159D : data <= 8'b00000000 ;
			15'h0000159E : data <= 8'b00000000 ;
			15'h0000159F : data <= 8'b00000000 ;
			15'h000015A0 : data <= 8'b00000000 ;
			15'h000015A1 : data <= 8'b00000000 ;
			15'h000015A2 : data <= 8'b00000000 ;
			15'h000015A3 : data <= 8'b00000000 ;
			15'h000015A4 : data <= 8'b00000000 ;
			15'h000015A5 : data <= 8'b00000000 ;
			15'h000015A6 : data <= 8'b00000000 ;
			15'h000015A7 : data <= 8'b00000000 ;
			15'h000015A8 : data <= 8'b00000000 ;
			15'h000015A9 : data <= 8'b00000000 ;
			15'h000015AA : data <= 8'b00000000 ;
			15'h000015AB : data <= 8'b00000000 ;
			15'h000015AC : data <= 8'b00000000 ;
			15'h000015AD : data <= 8'b00000000 ;
			15'h000015AE : data <= 8'b00000000 ;
			15'h000015AF : data <= 8'b00000000 ;
			15'h000015B0 : data <= 8'b00000000 ;
			15'h000015B1 : data <= 8'b00000000 ;
			15'h000015B2 : data <= 8'b00000000 ;
			15'h000015B3 : data <= 8'b00000000 ;
			15'h000015B4 : data <= 8'b00000000 ;
			15'h000015B5 : data <= 8'b00000000 ;
			15'h000015B6 : data <= 8'b00000000 ;
			15'h000015B7 : data <= 8'b00000000 ;
			15'h000015B8 : data <= 8'b00000000 ;
			15'h000015B9 : data <= 8'b00000000 ;
			15'h000015BA : data <= 8'b00000000 ;
			15'h000015BB : data <= 8'b00000000 ;
			15'h000015BC : data <= 8'b00000000 ;
			15'h000015BD : data <= 8'b00000000 ;
			15'h000015BE : data <= 8'b00000000 ;
			15'h000015BF : data <= 8'b00000000 ;
			15'h000015C0 : data <= 8'b00000000 ;
			15'h000015C1 : data <= 8'b00000000 ;
			15'h000015C2 : data <= 8'b00000000 ;
			15'h000015C3 : data <= 8'b00000000 ;
			15'h000015C4 : data <= 8'b00000000 ;
			15'h000015C5 : data <= 8'b00000000 ;
			15'h000015C6 : data <= 8'b00000000 ;
			15'h000015C7 : data <= 8'b00000000 ;
			15'h000015C8 : data <= 8'b00000000 ;
			15'h000015C9 : data <= 8'b00000000 ;
			15'h000015CA : data <= 8'b00000000 ;
			15'h000015CB : data <= 8'b00000000 ;
			15'h000015CC : data <= 8'b00000000 ;
			15'h000015CD : data <= 8'b00000000 ;
			15'h000015CE : data <= 8'b00000000 ;
			15'h000015CF : data <= 8'b00000000 ;
			15'h000015D0 : data <= 8'b00000000 ;
			15'h000015D1 : data <= 8'b00000000 ;
			15'h000015D2 : data <= 8'b00000000 ;
			15'h000015D3 : data <= 8'b00000000 ;
			15'h000015D4 : data <= 8'b00000000 ;
			15'h000015D5 : data <= 8'b00000000 ;
			15'h000015D6 : data <= 8'b00000000 ;
			15'h000015D7 : data <= 8'b00000000 ;
			15'h000015D8 : data <= 8'b00000000 ;
			15'h000015D9 : data <= 8'b00000000 ;
			15'h000015DA : data <= 8'b00000000 ;
			15'h000015DB : data <= 8'b00000000 ;
			15'h000015DC : data <= 8'b00000000 ;
			15'h000015DD : data <= 8'b00000000 ;
			15'h000015DE : data <= 8'b00000000 ;
			15'h000015DF : data <= 8'b00000000 ;
			15'h000015E0 : data <= 8'b00000000 ;
			15'h000015E1 : data <= 8'b00000000 ;
			15'h000015E2 : data <= 8'b00000000 ;
			15'h000015E3 : data <= 8'b00000000 ;
			15'h000015E4 : data <= 8'b00000000 ;
			15'h000015E5 : data <= 8'b00000000 ;
			15'h000015E6 : data <= 8'b00000000 ;
			15'h000015E7 : data <= 8'b00000000 ;
			15'h000015E8 : data <= 8'b00000000 ;
			15'h000015E9 : data <= 8'b00000000 ;
			15'h000015EA : data <= 8'b00000000 ;
			15'h000015EB : data <= 8'b00000000 ;
			15'h000015EC : data <= 8'b00000000 ;
			15'h000015ED : data <= 8'b00000000 ;
			15'h000015EE : data <= 8'b00000000 ;
			15'h000015EF : data <= 8'b00000000 ;
			15'h000015F0 : data <= 8'b00000000 ;
			15'h000015F1 : data <= 8'b00000000 ;
			15'h000015F2 : data <= 8'b00000000 ;
			15'h000015F3 : data <= 8'b00000000 ;
			15'h000015F4 : data <= 8'b00000000 ;
			15'h000015F5 : data <= 8'b00000000 ;
			15'h000015F6 : data <= 8'b00000000 ;
			15'h000015F7 : data <= 8'b00000000 ;
			15'h000015F8 : data <= 8'b00000000 ;
			15'h000015F9 : data <= 8'b00000000 ;
			15'h000015FA : data <= 8'b00000000 ;
			15'h000015FB : data <= 8'b00000000 ;
			15'h000015FC : data <= 8'b00000000 ;
			15'h000015FD : data <= 8'b00000000 ;
			15'h000015FE : data <= 8'b00000000 ;
			15'h000015FF : data <= 8'b00000000 ;
			15'h00001600 : data <= 8'b00000000 ;
			15'h00001601 : data <= 8'b00000000 ;
			15'h00001602 : data <= 8'b00000000 ;
			15'h00001603 : data <= 8'b00000000 ;
			15'h00001604 : data <= 8'b00000000 ;
			15'h00001605 : data <= 8'b00000000 ;
			15'h00001606 : data <= 8'b00000000 ;
			15'h00001607 : data <= 8'b00000000 ;
			15'h00001608 : data <= 8'b00000000 ;
			15'h00001609 : data <= 8'b00000000 ;
			15'h0000160A : data <= 8'b00000000 ;
			15'h0000160B : data <= 8'b00000000 ;
			15'h0000160C : data <= 8'b00000000 ;
			15'h0000160D : data <= 8'b00000000 ;
			15'h0000160E : data <= 8'b00000000 ;
			15'h0000160F : data <= 8'b00000000 ;
			15'h00001610 : data <= 8'b00000000 ;
			15'h00001611 : data <= 8'b00000000 ;
			15'h00001612 : data <= 8'b00000000 ;
			15'h00001613 : data <= 8'b00000000 ;
			15'h00001614 : data <= 8'b00000000 ;
			15'h00001615 : data <= 8'b00000000 ;
			15'h00001616 : data <= 8'b00000000 ;
			15'h00001617 : data <= 8'b00000000 ;
			15'h00001618 : data <= 8'b00000000 ;
			15'h00001619 : data <= 8'b00000000 ;
			15'h0000161A : data <= 8'b00000000 ;
			15'h0000161B : data <= 8'b00000000 ;
			15'h0000161C : data <= 8'b00000000 ;
			15'h0000161D : data <= 8'b00000000 ;
			15'h0000161E : data <= 8'b00000000 ;
			15'h0000161F : data <= 8'b00000000 ;
			15'h00001620 : data <= 8'b00000000 ;
			15'h00001621 : data <= 8'b00000000 ;
			15'h00001622 : data <= 8'b00000000 ;
			15'h00001623 : data <= 8'b00000000 ;
			15'h00001624 : data <= 8'b00000000 ;
			15'h00001625 : data <= 8'b00000000 ;
			15'h00001626 : data <= 8'b00000000 ;
			15'h00001627 : data <= 8'b00000000 ;
			15'h00001628 : data <= 8'b00000000 ;
			15'h00001629 : data <= 8'b00000000 ;
			15'h0000162A : data <= 8'b00000000 ;
			15'h0000162B : data <= 8'b00000000 ;
			15'h0000162C : data <= 8'b00000000 ;
			15'h0000162D : data <= 8'b00000000 ;
			15'h0000162E : data <= 8'b00000000 ;
			15'h0000162F : data <= 8'b00000000 ;
			15'h00001630 : data <= 8'b00000000 ;
			15'h00001631 : data <= 8'b00000000 ;
			15'h00001632 : data <= 8'b00000000 ;
			15'h00001633 : data <= 8'b00000000 ;
			15'h00001634 : data <= 8'b00000000 ;
			15'h00001635 : data <= 8'b00000000 ;
			15'h00001636 : data <= 8'b00000000 ;
			15'h00001637 : data <= 8'b00000000 ;
			15'h00001638 : data <= 8'b00000000 ;
			15'h00001639 : data <= 8'b00000000 ;
			15'h0000163A : data <= 8'b00000000 ;
			15'h0000163B : data <= 8'b00000000 ;
			15'h0000163C : data <= 8'b00000000 ;
			15'h0000163D : data <= 8'b00000000 ;
			15'h0000163E : data <= 8'b00000000 ;
			15'h0000163F : data <= 8'b00000000 ;
			15'h00001640 : data <= 8'b00000000 ;
			15'h00001641 : data <= 8'b00000000 ;
			15'h00001642 : data <= 8'b00000000 ;
			15'h00001643 : data <= 8'b00000000 ;
			15'h00001644 : data <= 8'b00000000 ;
			15'h00001645 : data <= 8'b00000000 ;
			15'h00001646 : data <= 8'b00000000 ;
			15'h00001647 : data <= 8'b00000000 ;
			15'h00001648 : data <= 8'b00000000 ;
			15'h00001649 : data <= 8'b00000000 ;
			15'h0000164A : data <= 8'b00000000 ;
			15'h0000164B : data <= 8'b00000000 ;
			15'h0000164C : data <= 8'b00000000 ;
			15'h0000164D : data <= 8'b00000000 ;
			15'h0000164E : data <= 8'b00000000 ;
			15'h0000164F : data <= 8'b00000000 ;
			15'h00001650 : data <= 8'b00000000 ;
			15'h00001651 : data <= 8'b00000000 ;
			15'h00001652 : data <= 8'b00000000 ;
			15'h00001653 : data <= 8'b00000000 ;
			15'h00001654 : data <= 8'b00000000 ;
			15'h00001655 : data <= 8'b00000000 ;
			15'h00001656 : data <= 8'b00000000 ;
			15'h00001657 : data <= 8'b00000000 ;
			15'h00001658 : data <= 8'b00000000 ;
			15'h00001659 : data <= 8'b00000000 ;
			15'h0000165A : data <= 8'b00000000 ;
			15'h0000165B : data <= 8'b00000000 ;
			15'h0000165C : data <= 8'b00000000 ;
			15'h0000165D : data <= 8'b00000000 ;
			15'h0000165E : data <= 8'b00000000 ;
			15'h0000165F : data <= 8'b00000000 ;
			15'h00001660 : data <= 8'b00000000 ;
			15'h00001661 : data <= 8'b00000000 ;
			15'h00001662 : data <= 8'b00000000 ;
			15'h00001663 : data <= 8'b00000000 ;
			15'h00001664 : data <= 8'b00000000 ;
			15'h00001665 : data <= 8'b00000000 ;
			15'h00001666 : data <= 8'b00000000 ;
			15'h00001667 : data <= 8'b00000000 ;
			15'h00001668 : data <= 8'b00000000 ;
			15'h00001669 : data <= 8'b00000000 ;
			15'h0000166A : data <= 8'b00000000 ;
			15'h0000166B : data <= 8'b00000000 ;
			15'h0000166C : data <= 8'b00000000 ;
			15'h0000166D : data <= 8'b00000000 ;
			15'h0000166E : data <= 8'b00000000 ;
			15'h0000166F : data <= 8'b00000000 ;
			15'h00001670 : data <= 8'b00000000 ;
			15'h00001671 : data <= 8'b00000000 ;
			15'h00001672 : data <= 8'b00000000 ;
			15'h00001673 : data <= 8'b00000000 ;
			15'h00001674 : data <= 8'b00000000 ;
			15'h00001675 : data <= 8'b00000000 ;
			15'h00001676 : data <= 8'b00000000 ;
			15'h00001677 : data <= 8'b00000000 ;
			15'h00001678 : data <= 8'b00000000 ;
			15'h00001679 : data <= 8'b00000000 ;
			15'h0000167A : data <= 8'b00000000 ;
			15'h0000167B : data <= 8'b00000000 ;
			15'h0000167C : data <= 8'b00000000 ;
			15'h0000167D : data <= 8'b00000000 ;
			15'h0000167E : data <= 8'b00000000 ;
			15'h0000167F : data <= 8'b00000000 ;
			15'h00001680 : data <= 8'b00000000 ;
			15'h00001681 : data <= 8'b00000000 ;
			15'h00001682 : data <= 8'b00000000 ;
			15'h00001683 : data <= 8'b00000000 ;
			15'h00001684 : data <= 8'b00000000 ;
			15'h00001685 : data <= 8'b00000000 ;
			15'h00001686 : data <= 8'b00000000 ;
			15'h00001687 : data <= 8'b00000000 ;
			15'h00001688 : data <= 8'b00000000 ;
			15'h00001689 : data <= 8'b00000000 ;
			15'h0000168A : data <= 8'b00000000 ;
			15'h0000168B : data <= 8'b00000000 ;
			15'h0000168C : data <= 8'b00000000 ;
			15'h0000168D : data <= 8'b00000000 ;
			15'h0000168E : data <= 8'b00000000 ;
			15'h0000168F : data <= 8'b00000000 ;
			15'h00001690 : data <= 8'b00000000 ;
			15'h00001691 : data <= 8'b00000000 ;
			15'h00001692 : data <= 8'b00000000 ;
			15'h00001693 : data <= 8'b00000000 ;
			15'h00001694 : data <= 8'b00000000 ;
			15'h00001695 : data <= 8'b00000000 ;
			15'h00001696 : data <= 8'b00000000 ;
			15'h00001697 : data <= 8'b00000000 ;
			15'h00001698 : data <= 8'b00000000 ;
			15'h00001699 : data <= 8'b00000000 ;
			15'h0000169A : data <= 8'b00000000 ;
			15'h0000169B : data <= 8'b00000000 ;
			15'h0000169C : data <= 8'b00000000 ;
			15'h0000169D : data <= 8'b00000000 ;
			15'h0000169E : data <= 8'b00000000 ;
			15'h0000169F : data <= 8'b00000000 ;
			15'h000016A0 : data <= 8'b00000000 ;
			15'h000016A1 : data <= 8'b00000000 ;
			15'h000016A2 : data <= 8'b00000000 ;
			15'h000016A3 : data <= 8'b00000000 ;
			15'h000016A4 : data <= 8'b00000000 ;
			15'h000016A5 : data <= 8'b00000000 ;
			15'h000016A6 : data <= 8'b00000000 ;
			15'h000016A7 : data <= 8'b00000000 ;
			15'h000016A8 : data <= 8'b00000000 ;
			15'h000016A9 : data <= 8'b00000000 ;
			15'h000016AA : data <= 8'b00000000 ;
			15'h000016AB : data <= 8'b00000000 ;
			15'h000016AC : data <= 8'b00000000 ;
			15'h000016AD : data <= 8'b00000000 ;
			15'h000016AE : data <= 8'b00000000 ;
			15'h000016AF : data <= 8'b00000000 ;
			15'h000016B0 : data <= 8'b00000000 ;
			15'h000016B1 : data <= 8'b00000000 ;
			15'h000016B2 : data <= 8'b00000000 ;
			15'h000016B3 : data <= 8'b00000000 ;
			15'h000016B4 : data <= 8'b00000000 ;
			15'h000016B5 : data <= 8'b00000000 ;
			15'h000016B6 : data <= 8'b00000000 ;
			15'h000016B7 : data <= 8'b00000000 ;
			15'h000016B8 : data <= 8'b00000000 ;
			15'h000016B9 : data <= 8'b00000000 ;
			15'h000016BA : data <= 8'b00000000 ;
			15'h000016BB : data <= 8'b00000000 ;
			15'h000016BC : data <= 8'b00000000 ;
			15'h000016BD : data <= 8'b00000000 ;
			15'h000016BE : data <= 8'b00000000 ;
			15'h000016BF : data <= 8'b00000000 ;
			15'h000016C0 : data <= 8'b00000000 ;
			15'h000016C1 : data <= 8'b00000000 ;
			15'h000016C2 : data <= 8'b00000000 ;
			15'h000016C3 : data <= 8'b00000000 ;
			15'h000016C4 : data <= 8'b00000000 ;
			15'h000016C5 : data <= 8'b00000000 ;
			15'h000016C6 : data <= 8'b00000000 ;
			15'h000016C7 : data <= 8'b00000000 ;
			15'h000016C8 : data <= 8'b00000000 ;
			15'h000016C9 : data <= 8'b00000000 ;
			15'h000016CA : data <= 8'b00000000 ;
			15'h000016CB : data <= 8'b00000000 ;
			15'h000016CC : data <= 8'b00000000 ;
			15'h000016CD : data <= 8'b00000000 ;
			15'h000016CE : data <= 8'b00000000 ;
			15'h000016CF : data <= 8'b00000000 ;
			15'h000016D0 : data <= 8'b00000000 ;
			15'h000016D1 : data <= 8'b00000000 ;
			15'h000016D2 : data <= 8'b00000000 ;
			15'h000016D3 : data <= 8'b00000000 ;
			15'h000016D4 : data <= 8'b00000000 ;
			15'h000016D5 : data <= 8'b00000000 ;
			15'h000016D6 : data <= 8'b00000000 ;
			15'h000016D7 : data <= 8'b00000000 ;
			15'h000016D8 : data <= 8'b00000000 ;
			15'h000016D9 : data <= 8'b00000000 ;
			15'h000016DA : data <= 8'b00000000 ;
			15'h000016DB : data <= 8'b00000000 ;
			15'h000016DC : data <= 8'b00000000 ;
			15'h000016DD : data <= 8'b00000000 ;
			15'h000016DE : data <= 8'b00000000 ;
			15'h000016DF : data <= 8'b00000000 ;
			15'h000016E0 : data <= 8'b00000000 ;
			15'h000016E1 : data <= 8'b00000000 ;
			15'h000016E2 : data <= 8'b00000000 ;
			15'h000016E3 : data <= 8'b00000000 ;
			15'h000016E4 : data <= 8'b00000000 ;
			15'h000016E5 : data <= 8'b00000000 ;
			15'h000016E6 : data <= 8'b00000000 ;
			15'h000016E7 : data <= 8'b00000000 ;
			15'h000016E8 : data <= 8'b00000000 ;
			15'h000016E9 : data <= 8'b00000000 ;
			15'h000016EA : data <= 8'b00000000 ;
			15'h000016EB : data <= 8'b00000000 ;
			15'h000016EC : data <= 8'b00000000 ;
			15'h000016ED : data <= 8'b00000000 ;
			15'h000016EE : data <= 8'b00000000 ;
			15'h000016EF : data <= 8'b00000000 ;
			15'h000016F0 : data <= 8'b00000000 ;
			15'h000016F1 : data <= 8'b00000000 ;
			15'h000016F2 : data <= 8'b00000000 ;
			15'h000016F3 : data <= 8'b00000000 ;
			15'h000016F4 : data <= 8'b00000000 ;
			15'h000016F5 : data <= 8'b00000000 ;
			15'h000016F6 : data <= 8'b00000000 ;
			15'h000016F7 : data <= 8'b00000000 ;
			15'h000016F8 : data <= 8'b00000000 ;
			15'h000016F9 : data <= 8'b00000000 ;
			15'h000016FA : data <= 8'b00000000 ;
			15'h000016FB : data <= 8'b00000000 ;
			15'h000016FC : data <= 8'b00000000 ;
			15'h000016FD : data <= 8'b00000000 ;
			15'h000016FE : data <= 8'b00000000 ;
			15'h000016FF : data <= 8'b00000000 ;
			15'h00001700 : data <= 8'b00000000 ;
			15'h00001701 : data <= 8'b00000000 ;
			15'h00001702 : data <= 8'b00000000 ;
			15'h00001703 : data <= 8'b00000000 ;
			15'h00001704 : data <= 8'b00000000 ;
			15'h00001705 : data <= 8'b00000000 ;
			15'h00001706 : data <= 8'b00000000 ;
			15'h00001707 : data <= 8'b00000000 ;
			15'h00001708 : data <= 8'b00000000 ;
			15'h00001709 : data <= 8'b00000000 ;
			15'h0000170A : data <= 8'b00000000 ;
			15'h0000170B : data <= 8'b00000000 ;
			15'h0000170C : data <= 8'b00000000 ;
			15'h0000170D : data <= 8'b00000000 ;
			15'h0000170E : data <= 8'b00000000 ;
			15'h0000170F : data <= 8'b00000000 ;
			15'h00001710 : data <= 8'b00000000 ;
			15'h00001711 : data <= 8'b00000000 ;
			15'h00001712 : data <= 8'b00000000 ;
			15'h00001713 : data <= 8'b00000000 ;
			15'h00001714 : data <= 8'b00000000 ;
			15'h00001715 : data <= 8'b00000000 ;
			15'h00001716 : data <= 8'b00000000 ;
			15'h00001717 : data <= 8'b00000000 ;
			15'h00001718 : data <= 8'b00000000 ;
			15'h00001719 : data <= 8'b00000000 ;
			15'h0000171A : data <= 8'b00000000 ;
			15'h0000171B : data <= 8'b00000000 ;
			15'h0000171C : data <= 8'b00000000 ;
			15'h0000171D : data <= 8'b00000000 ;
			15'h0000171E : data <= 8'b00000000 ;
			15'h0000171F : data <= 8'b00000000 ;
			15'h00001720 : data <= 8'b00000000 ;
			15'h00001721 : data <= 8'b00000000 ;
			15'h00001722 : data <= 8'b00000000 ;
			15'h00001723 : data <= 8'b00000000 ;
			15'h00001724 : data <= 8'b00000000 ;
			15'h00001725 : data <= 8'b00000000 ;
			15'h00001726 : data <= 8'b00000000 ;
			15'h00001727 : data <= 8'b00000000 ;
			15'h00001728 : data <= 8'b00000000 ;
			15'h00001729 : data <= 8'b00000000 ;
			15'h0000172A : data <= 8'b00000000 ;
			15'h0000172B : data <= 8'b00000000 ;
			15'h0000172C : data <= 8'b00000000 ;
			15'h0000172D : data <= 8'b00000000 ;
			15'h0000172E : data <= 8'b00000000 ;
			15'h0000172F : data <= 8'b00000000 ;
			15'h00001730 : data <= 8'b00000000 ;
			15'h00001731 : data <= 8'b00000000 ;
			15'h00001732 : data <= 8'b00000000 ;
			15'h00001733 : data <= 8'b00000000 ;
			15'h00001734 : data <= 8'b00000000 ;
			15'h00001735 : data <= 8'b00000000 ;
			15'h00001736 : data <= 8'b00000000 ;
			15'h00001737 : data <= 8'b00000000 ;
			15'h00001738 : data <= 8'b00000000 ;
			15'h00001739 : data <= 8'b00000000 ;
			15'h0000173A : data <= 8'b00000000 ;
			15'h0000173B : data <= 8'b00000000 ;
			15'h0000173C : data <= 8'b00000000 ;
			15'h0000173D : data <= 8'b00000000 ;
			15'h0000173E : data <= 8'b00000000 ;
			15'h0000173F : data <= 8'b00000000 ;
			15'h00001740 : data <= 8'b00000000 ;
			15'h00001741 : data <= 8'b00000000 ;
			15'h00001742 : data <= 8'b00000000 ;
			15'h00001743 : data <= 8'b00000000 ;
			15'h00001744 : data <= 8'b00000000 ;
			15'h00001745 : data <= 8'b00000000 ;
			15'h00001746 : data <= 8'b00000000 ;
			15'h00001747 : data <= 8'b00000000 ;
			15'h00001748 : data <= 8'b00000000 ;
			15'h00001749 : data <= 8'b00000000 ;
			15'h0000174A : data <= 8'b00000000 ;
			15'h0000174B : data <= 8'b00000000 ;
			15'h0000174C : data <= 8'b00000000 ;
			15'h0000174D : data <= 8'b00000000 ;
			15'h0000174E : data <= 8'b00000000 ;
			15'h0000174F : data <= 8'b00000000 ;
			15'h00001750 : data <= 8'b00000000 ;
			15'h00001751 : data <= 8'b00000000 ;
			15'h00001752 : data <= 8'b00000000 ;
			15'h00001753 : data <= 8'b00000000 ;
			15'h00001754 : data <= 8'b00000000 ;
			15'h00001755 : data <= 8'b00000000 ;
			15'h00001756 : data <= 8'b00000000 ;
			15'h00001757 : data <= 8'b00000000 ;
			15'h00001758 : data <= 8'b00000000 ;
			15'h00001759 : data <= 8'b00000000 ;
			15'h0000175A : data <= 8'b00000000 ;
			15'h0000175B : data <= 8'b00000000 ;
			15'h0000175C : data <= 8'b00000000 ;
			15'h0000175D : data <= 8'b00000000 ;
			15'h0000175E : data <= 8'b00000000 ;
			15'h0000175F : data <= 8'b00000000 ;
			15'h00001760 : data <= 8'b00000000 ;
			15'h00001761 : data <= 8'b00000000 ;
			15'h00001762 : data <= 8'b00000000 ;
			15'h00001763 : data <= 8'b00000000 ;
			15'h00001764 : data <= 8'b00000000 ;
			15'h00001765 : data <= 8'b00000000 ;
			15'h00001766 : data <= 8'b00000000 ;
			15'h00001767 : data <= 8'b00000000 ;
			15'h00001768 : data <= 8'b00000000 ;
			15'h00001769 : data <= 8'b00000000 ;
			15'h0000176A : data <= 8'b00000000 ;
			15'h0000176B : data <= 8'b00000000 ;
			15'h0000176C : data <= 8'b00000000 ;
			15'h0000176D : data <= 8'b00000000 ;
			15'h0000176E : data <= 8'b00000000 ;
			15'h0000176F : data <= 8'b00000000 ;
			15'h00001770 : data <= 8'b00000000 ;
			15'h00001771 : data <= 8'b00000000 ;
			15'h00001772 : data <= 8'b00000000 ;
			15'h00001773 : data <= 8'b00000000 ;
			15'h00001774 : data <= 8'b00000000 ;
			15'h00001775 : data <= 8'b00000000 ;
			15'h00001776 : data <= 8'b00000000 ;
			15'h00001777 : data <= 8'b00000000 ;
			15'h00001778 : data <= 8'b00000000 ;
			15'h00001779 : data <= 8'b00000000 ;
			15'h0000177A : data <= 8'b00000000 ;
			15'h0000177B : data <= 8'b00000000 ;
			15'h0000177C : data <= 8'b00000000 ;
			15'h0000177D : data <= 8'b00000000 ;
			15'h0000177E : data <= 8'b00000000 ;
			15'h0000177F : data <= 8'b00000000 ;
			15'h00001780 : data <= 8'b00000000 ;
			15'h00001781 : data <= 8'b00000000 ;
			15'h00001782 : data <= 8'b00000000 ;
			15'h00001783 : data <= 8'b00000000 ;
			15'h00001784 : data <= 8'b00000000 ;
			15'h00001785 : data <= 8'b00000000 ;
			15'h00001786 : data <= 8'b00000000 ;
			15'h00001787 : data <= 8'b00000000 ;
			15'h00001788 : data <= 8'b00000000 ;
			15'h00001789 : data <= 8'b00000000 ;
			15'h0000178A : data <= 8'b00000000 ;
			15'h0000178B : data <= 8'b00000000 ;
			15'h0000178C : data <= 8'b00000000 ;
			15'h0000178D : data <= 8'b00000000 ;
			15'h0000178E : data <= 8'b00000000 ;
			15'h0000178F : data <= 8'b00000000 ;
			15'h00001790 : data <= 8'b00000000 ;
			15'h00001791 : data <= 8'b00000000 ;
			15'h00001792 : data <= 8'b00000000 ;
			15'h00001793 : data <= 8'b00000000 ;
			15'h00001794 : data <= 8'b00000000 ;
			15'h00001795 : data <= 8'b00000000 ;
			15'h00001796 : data <= 8'b00000000 ;
			15'h00001797 : data <= 8'b00000000 ;
			15'h00001798 : data <= 8'b00000000 ;
			15'h00001799 : data <= 8'b00000000 ;
			15'h0000179A : data <= 8'b00000000 ;
			15'h0000179B : data <= 8'b00000000 ;
			15'h0000179C : data <= 8'b00000000 ;
			15'h0000179D : data <= 8'b00000000 ;
			15'h0000179E : data <= 8'b00000000 ;
			15'h0000179F : data <= 8'b00000000 ;
			15'h000017A0 : data <= 8'b00000000 ;
			15'h000017A1 : data <= 8'b00000000 ;
			15'h000017A2 : data <= 8'b00000000 ;
			15'h000017A3 : data <= 8'b00000000 ;
			15'h000017A4 : data <= 8'b00000000 ;
			15'h000017A5 : data <= 8'b00000000 ;
			15'h000017A6 : data <= 8'b00000000 ;
			15'h000017A7 : data <= 8'b00000000 ;
			15'h000017A8 : data <= 8'b00000000 ;
			15'h000017A9 : data <= 8'b00000000 ;
			15'h000017AA : data <= 8'b00000000 ;
			15'h000017AB : data <= 8'b00000000 ;
			15'h000017AC : data <= 8'b00000000 ;
			15'h000017AD : data <= 8'b00000000 ;
			15'h000017AE : data <= 8'b00000000 ;
			15'h000017AF : data <= 8'b00000000 ;
			15'h000017B0 : data <= 8'b00000000 ;
			15'h000017B1 : data <= 8'b00000000 ;
			15'h000017B2 : data <= 8'b00000000 ;
			15'h000017B3 : data <= 8'b00000000 ;
			15'h000017B4 : data <= 8'b00000000 ;
			15'h000017B5 : data <= 8'b00000000 ;
			15'h000017B6 : data <= 8'b00000000 ;
			15'h000017B7 : data <= 8'b00000000 ;
			15'h000017B8 : data <= 8'b00000000 ;
			15'h000017B9 : data <= 8'b00000000 ;
			15'h000017BA : data <= 8'b00000000 ;
			15'h000017BB : data <= 8'b00000000 ;
			15'h000017BC : data <= 8'b00000000 ;
			15'h000017BD : data <= 8'b00000000 ;
			15'h000017BE : data <= 8'b00000000 ;
			15'h000017BF : data <= 8'b00000000 ;
			15'h000017C0 : data <= 8'b00000000 ;
			15'h000017C1 : data <= 8'b00000000 ;
			15'h000017C2 : data <= 8'b00000000 ;
			15'h000017C3 : data <= 8'b00000000 ;
			15'h000017C4 : data <= 8'b00000000 ;
			15'h000017C5 : data <= 8'b00000000 ;
			15'h000017C6 : data <= 8'b00000000 ;
			15'h000017C7 : data <= 8'b00000000 ;
			15'h000017C8 : data <= 8'b00000000 ;
			15'h000017C9 : data <= 8'b00000000 ;
			15'h000017CA : data <= 8'b00000000 ;
			15'h000017CB : data <= 8'b00000000 ;
			15'h000017CC : data <= 8'b00000000 ;
			15'h000017CD : data <= 8'b00000000 ;
			15'h000017CE : data <= 8'b00000000 ;
			15'h000017CF : data <= 8'b00000000 ;
			15'h000017D0 : data <= 8'b00000000 ;
			15'h000017D1 : data <= 8'b00000000 ;
			15'h000017D2 : data <= 8'b00000000 ;
			15'h000017D3 : data <= 8'b00000000 ;
			15'h000017D4 : data <= 8'b00000000 ;
			15'h000017D5 : data <= 8'b00000000 ;
			15'h000017D6 : data <= 8'b00000000 ;
			15'h000017D7 : data <= 8'b00000000 ;
			15'h000017D8 : data <= 8'b00000000 ;
			15'h000017D9 : data <= 8'b00000000 ;
			15'h000017DA : data <= 8'b00000000 ;
			15'h000017DB : data <= 8'b00000000 ;
			15'h000017DC : data <= 8'b00000000 ;
			15'h000017DD : data <= 8'b00000000 ;
			15'h000017DE : data <= 8'b00000000 ;
			15'h000017DF : data <= 8'b00000000 ;
			15'h000017E0 : data <= 8'b00000000 ;
			15'h000017E1 : data <= 8'b00000000 ;
			15'h000017E2 : data <= 8'b00000000 ;
			15'h000017E3 : data <= 8'b00000000 ;
			15'h000017E4 : data <= 8'b00000000 ;
			15'h000017E5 : data <= 8'b00000000 ;
			15'h000017E6 : data <= 8'b00000000 ;
			15'h000017E7 : data <= 8'b00000000 ;
			15'h000017E8 : data <= 8'b00000000 ;
			15'h000017E9 : data <= 8'b00000000 ;
			15'h000017EA : data <= 8'b00000000 ;
			15'h000017EB : data <= 8'b00000000 ;
			15'h000017EC : data <= 8'b00000000 ;
			15'h000017ED : data <= 8'b00000000 ;
			15'h000017EE : data <= 8'b00000000 ;
			15'h000017EF : data <= 8'b00000000 ;
			15'h000017F0 : data <= 8'b00000000 ;
			15'h000017F1 : data <= 8'b00000000 ;
			15'h000017F2 : data <= 8'b00000000 ;
			15'h000017F3 : data <= 8'b00000000 ;
			15'h000017F4 : data <= 8'b00000000 ;
			15'h000017F5 : data <= 8'b00000000 ;
			15'h000017F6 : data <= 8'b00000000 ;
			15'h000017F7 : data <= 8'b00000000 ;
			15'h000017F8 : data <= 8'b00000000 ;
			15'h000017F9 : data <= 8'b00000000 ;
			15'h000017FA : data <= 8'b00000000 ;
			15'h000017FB : data <= 8'b00000000 ;
			15'h000017FC : data <= 8'b00000000 ;
			15'h000017FD : data <= 8'b00000000 ;
			15'h000017FE : data <= 8'b00000000 ;
			15'h000017FF : data <= 8'b00000000 ;
			15'h00001800 : data <= 8'b00000000 ;
			15'h00001801 : data <= 8'b00000000 ;
			15'h00001802 : data <= 8'b00000000 ;
			15'h00001803 : data <= 8'b00000000 ;
			15'h00001804 : data <= 8'b00000000 ;
			15'h00001805 : data <= 8'b00000000 ;
			15'h00001806 : data <= 8'b00000000 ;
			15'h00001807 : data <= 8'b00000000 ;
			15'h00001808 : data <= 8'b00000000 ;
			15'h00001809 : data <= 8'b00000000 ;
			15'h0000180A : data <= 8'b00000000 ;
			15'h0000180B : data <= 8'b00000000 ;
			15'h0000180C : data <= 8'b00000000 ;
			15'h0000180D : data <= 8'b00000000 ;
			15'h0000180E : data <= 8'b00000000 ;
			15'h0000180F : data <= 8'b00000000 ;
			15'h00001810 : data <= 8'b00000000 ;
			15'h00001811 : data <= 8'b00000000 ;
			15'h00001812 : data <= 8'b00000000 ;
			15'h00001813 : data <= 8'b00000000 ;
			15'h00001814 : data <= 8'b00000000 ;
			15'h00001815 : data <= 8'b00000000 ;
			15'h00001816 : data <= 8'b00000000 ;
			15'h00001817 : data <= 8'b00000000 ;
			15'h00001818 : data <= 8'b00000000 ;
			15'h00001819 : data <= 8'b00000000 ;
			15'h0000181A : data <= 8'b00000000 ;
			15'h0000181B : data <= 8'b00000000 ;
			15'h0000181C : data <= 8'b00000000 ;
			15'h0000181D : data <= 8'b00000000 ;
			15'h0000181E : data <= 8'b00000000 ;
			15'h0000181F : data <= 8'b00000000 ;
			15'h00001820 : data <= 8'b00000000 ;
			15'h00001821 : data <= 8'b00000000 ;
			15'h00001822 : data <= 8'b00000000 ;
			15'h00001823 : data <= 8'b00000000 ;
			15'h00001824 : data <= 8'b00000000 ;
			15'h00001825 : data <= 8'b00000000 ;
			15'h00001826 : data <= 8'b00000000 ;
			15'h00001827 : data <= 8'b00000000 ;
			15'h00001828 : data <= 8'b00000000 ;
			15'h00001829 : data <= 8'b00000000 ;
			15'h0000182A : data <= 8'b00000000 ;
			15'h0000182B : data <= 8'b00000000 ;
			15'h0000182C : data <= 8'b00000000 ;
			15'h0000182D : data <= 8'b00000000 ;
			15'h0000182E : data <= 8'b00000000 ;
			15'h0000182F : data <= 8'b00000000 ;
			15'h00001830 : data <= 8'b00000000 ;
			15'h00001831 : data <= 8'b00000000 ;
			15'h00001832 : data <= 8'b00000000 ;
			15'h00001833 : data <= 8'b00000000 ;
			15'h00001834 : data <= 8'b00000000 ;
			15'h00001835 : data <= 8'b00000000 ;
			15'h00001836 : data <= 8'b00000000 ;
			15'h00001837 : data <= 8'b00000000 ;
			15'h00001838 : data <= 8'b00000000 ;
			15'h00001839 : data <= 8'b00000000 ;
			15'h0000183A : data <= 8'b00000000 ;
			15'h0000183B : data <= 8'b00000000 ;
			15'h0000183C : data <= 8'b00000000 ;
			15'h0000183D : data <= 8'b00000000 ;
			15'h0000183E : data <= 8'b00000000 ;
			15'h0000183F : data <= 8'b00000000 ;
			15'h00001840 : data <= 8'b00000000 ;
			15'h00001841 : data <= 8'b00000000 ;
			15'h00001842 : data <= 8'b00000000 ;
			15'h00001843 : data <= 8'b00000000 ;
			15'h00001844 : data <= 8'b00000000 ;
			15'h00001845 : data <= 8'b00000000 ;
			15'h00001846 : data <= 8'b00000000 ;
			15'h00001847 : data <= 8'b00000000 ;
			15'h00001848 : data <= 8'b00000000 ;
			15'h00001849 : data <= 8'b00000000 ;
			15'h0000184A : data <= 8'b00000000 ;
			15'h0000184B : data <= 8'b00000000 ;
			15'h0000184C : data <= 8'b00000000 ;
			15'h0000184D : data <= 8'b00000000 ;
			15'h0000184E : data <= 8'b00000000 ;
			15'h0000184F : data <= 8'b00000000 ;
			15'h00001850 : data <= 8'b00000000 ;
			15'h00001851 : data <= 8'b00000000 ;
			15'h00001852 : data <= 8'b00000000 ;
			15'h00001853 : data <= 8'b00000000 ;
			15'h00001854 : data <= 8'b00000000 ;
			15'h00001855 : data <= 8'b00000000 ;
			15'h00001856 : data <= 8'b00000000 ;
			15'h00001857 : data <= 8'b00000000 ;
			15'h00001858 : data <= 8'b00000000 ;
			15'h00001859 : data <= 8'b00000000 ;
			15'h0000185A : data <= 8'b00000000 ;
			15'h0000185B : data <= 8'b00000000 ;
			15'h0000185C : data <= 8'b00000000 ;
			15'h0000185D : data <= 8'b00000000 ;
			15'h0000185E : data <= 8'b00000000 ;
			15'h0000185F : data <= 8'b00000000 ;
			15'h00001860 : data <= 8'b00000000 ;
			15'h00001861 : data <= 8'b00000000 ;
			15'h00001862 : data <= 8'b00000000 ;
			15'h00001863 : data <= 8'b00000000 ;
			15'h00001864 : data <= 8'b00000000 ;
			15'h00001865 : data <= 8'b00000000 ;
			15'h00001866 : data <= 8'b00000000 ;
			15'h00001867 : data <= 8'b00000000 ;
			15'h00001868 : data <= 8'b00000000 ;
			15'h00001869 : data <= 8'b00000000 ;
			15'h0000186A : data <= 8'b00000000 ;
			15'h0000186B : data <= 8'b00000000 ;
			15'h0000186C : data <= 8'b00000000 ;
			15'h0000186D : data <= 8'b00000000 ;
			15'h0000186E : data <= 8'b00000000 ;
			15'h0000186F : data <= 8'b00000000 ;
			15'h00001870 : data <= 8'b00000000 ;
			15'h00001871 : data <= 8'b00000000 ;
			15'h00001872 : data <= 8'b00000000 ;
			15'h00001873 : data <= 8'b00000000 ;
			15'h00001874 : data <= 8'b00000000 ;
			15'h00001875 : data <= 8'b00000000 ;
			15'h00001876 : data <= 8'b00000000 ;
			15'h00001877 : data <= 8'b00000000 ;
			15'h00001878 : data <= 8'b00000000 ;
			15'h00001879 : data <= 8'b00000000 ;
			15'h0000187A : data <= 8'b00000000 ;
			15'h0000187B : data <= 8'b00000000 ;
			15'h0000187C : data <= 8'b00000000 ;
			15'h0000187D : data <= 8'b00000000 ;
			15'h0000187E : data <= 8'b00000000 ;
			15'h0000187F : data <= 8'b00000000 ;
			15'h00001880 : data <= 8'b00000000 ;
			15'h00001881 : data <= 8'b00000000 ;
			15'h00001882 : data <= 8'b00000000 ;
			15'h00001883 : data <= 8'b00000000 ;
			15'h00001884 : data <= 8'b00000000 ;
			15'h00001885 : data <= 8'b00000000 ;
			15'h00001886 : data <= 8'b00000000 ;
			15'h00001887 : data <= 8'b00000000 ;
			15'h00001888 : data <= 8'b00000000 ;
			15'h00001889 : data <= 8'b00000000 ;
			15'h0000188A : data <= 8'b00000000 ;
			15'h0000188B : data <= 8'b00000000 ;
			15'h0000188C : data <= 8'b00000000 ;
			15'h0000188D : data <= 8'b00000000 ;
			15'h0000188E : data <= 8'b00000000 ;
			15'h0000188F : data <= 8'b00000000 ;
			15'h00001890 : data <= 8'b00000000 ;
			15'h00001891 : data <= 8'b00000000 ;
			15'h00001892 : data <= 8'b00000000 ;
			15'h00001893 : data <= 8'b00000000 ;
			15'h00001894 : data <= 8'b00000000 ;
			15'h00001895 : data <= 8'b00000000 ;
			15'h00001896 : data <= 8'b00000000 ;
			15'h00001897 : data <= 8'b00000000 ;
			15'h00001898 : data <= 8'b00000000 ;
			15'h00001899 : data <= 8'b00000000 ;
			15'h0000189A : data <= 8'b00000000 ;
			15'h0000189B : data <= 8'b00000000 ;
			15'h0000189C : data <= 8'b00000000 ;
			15'h0000189D : data <= 8'b00000000 ;
			15'h0000189E : data <= 8'b00000000 ;
			15'h0000189F : data <= 8'b00000000 ;
			15'h000018A0 : data <= 8'b00000000 ;
			15'h000018A1 : data <= 8'b00000000 ;
			15'h000018A2 : data <= 8'b00000000 ;
			15'h000018A3 : data <= 8'b00000000 ;
			15'h000018A4 : data <= 8'b00000000 ;
			15'h000018A5 : data <= 8'b00000000 ;
			15'h000018A6 : data <= 8'b00000000 ;
			15'h000018A7 : data <= 8'b00000000 ;
			15'h000018A8 : data <= 8'b00000000 ;
			15'h000018A9 : data <= 8'b00000000 ;
			15'h000018AA : data <= 8'b00000000 ;
			15'h000018AB : data <= 8'b00000000 ;
			15'h000018AC : data <= 8'b00000000 ;
			15'h000018AD : data <= 8'b00000000 ;
			15'h000018AE : data <= 8'b00000000 ;
			15'h000018AF : data <= 8'b00000000 ;
			15'h000018B0 : data <= 8'b00000000 ;
			15'h000018B1 : data <= 8'b00000000 ;
			15'h000018B2 : data <= 8'b00000000 ;
			15'h000018B3 : data <= 8'b00000000 ;
			15'h000018B4 : data <= 8'b00000000 ;
			15'h000018B5 : data <= 8'b00000000 ;
			15'h000018B6 : data <= 8'b00000000 ;
			15'h000018B7 : data <= 8'b00000000 ;
			15'h000018B8 : data <= 8'b00000000 ;
			15'h000018B9 : data <= 8'b00000000 ;
			15'h000018BA : data <= 8'b00000000 ;
			15'h000018BB : data <= 8'b00000000 ;
			15'h000018BC : data <= 8'b00000000 ;
			15'h000018BD : data <= 8'b00000000 ;
			15'h000018BE : data <= 8'b00000000 ;
			15'h000018BF : data <= 8'b00000000 ;
			15'h000018C0 : data <= 8'b00000000 ;
			15'h000018C1 : data <= 8'b00000000 ;
			15'h000018C2 : data <= 8'b00000000 ;
			15'h000018C3 : data <= 8'b00000000 ;
			15'h000018C4 : data <= 8'b00000000 ;
			15'h000018C5 : data <= 8'b00000000 ;
			15'h000018C6 : data <= 8'b00000000 ;
			15'h000018C7 : data <= 8'b00000000 ;
			15'h000018C8 : data <= 8'b00000000 ;
			15'h000018C9 : data <= 8'b00000000 ;
			15'h000018CA : data <= 8'b00000000 ;
			15'h000018CB : data <= 8'b00000000 ;
			15'h000018CC : data <= 8'b00000000 ;
			15'h000018CD : data <= 8'b00000000 ;
			15'h000018CE : data <= 8'b00000000 ;
			15'h000018CF : data <= 8'b00000000 ;
			15'h000018D0 : data <= 8'b00000000 ;
			15'h000018D1 : data <= 8'b00000000 ;
			15'h000018D2 : data <= 8'b00000000 ;
			15'h000018D3 : data <= 8'b00000000 ;
			15'h000018D4 : data <= 8'b00000000 ;
			15'h000018D5 : data <= 8'b00000000 ;
			15'h000018D6 : data <= 8'b00000000 ;
			15'h000018D7 : data <= 8'b00000000 ;
			15'h000018D8 : data <= 8'b00000000 ;
			15'h000018D9 : data <= 8'b00000000 ;
			15'h000018DA : data <= 8'b00000000 ;
			15'h000018DB : data <= 8'b00000000 ;
			15'h000018DC : data <= 8'b00000000 ;
			15'h000018DD : data <= 8'b00000000 ;
			15'h000018DE : data <= 8'b00000000 ;
			15'h000018DF : data <= 8'b00000000 ;
			15'h000018E0 : data <= 8'b00000000 ;
			15'h000018E1 : data <= 8'b00000000 ;
			15'h000018E2 : data <= 8'b00000000 ;
			15'h000018E3 : data <= 8'b00000000 ;
			15'h000018E4 : data <= 8'b00000000 ;
			15'h000018E5 : data <= 8'b00000000 ;
			15'h000018E6 : data <= 8'b00000000 ;
			15'h000018E7 : data <= 8'b00000000 ;
			15'h000018E8 : data <= 8'b00000000 ;
			15'h000018E9 : data <= 8'b00000000 ;
			15'h000018EA : data <= 8'b00000000 ;
			15'h000018EB : data <= 8'b00000000 ;
			15'h000018EC : data <= 8'b00000000 ;
			15'h000018ED : data <= 8'b00000000 ;
			15'h000018EE : data <= 8'b00000000 ;
			15'h000018EF : data <= 8'b00000000 ;
			15'h000018F0 : data <= 8'b00000000 ;
			15'h000018F1 : data <= 8'b00000000 ;
			15'h000018F2 : data <= 8'b00000000 ;
			15'h000018F3 : data <= 8'b00000000 ;
			15'h000018F4 : data <= 8'b00000000 ;
			15'h000018F5 : data <= 8'b00000000 ;
			15'h000018F6 : data <= 8'b00000000 ;
			15'h000018F7 : data <= 8'b00000000 ;
			15'h000018F8 : data <= 8'b00000000 ;
			15'h000018F9 : data <= 8'b00000000 ;
			15'h000018FA : data <= 8'b00000000 ;
			15'h000018FB : data <= 8'b00000000 ;
			15'h000018FC : data <= 8'b00000000 ;
			15'h000018FD : data <= 8'b00000000 ;
			15'h000018FE : data <= 8'b00000000 ;
			15'h000018FF : data <= 8'b00000000 ;
			15'h00001900 : data <= 8'b00000000 ;
			15'h00001901 : data <= 8'b00000000 ;
			15'h00001902 : data <= 8'b00000000 ;
			15'h00001903 : data <= 8'b00000000 ;
			15'h00001904 : data <= 8'b00000000 ;
			15'h00001905 : data <= 8'b00000000 ;
			15'h00001906 : data <= 8'b00000000 ;
			15'h00001907 : data <= 8'b00000000 ;
			15'h00001908 : data <= 8'b00000000 ;
			15'h00001909 : data <= 8'b00000000 ;
			15'h0000190A : data <= 8'b00000000 ;
			15'h0000190B : data <= 8'b00000000 ;
			15'h0000190C : data <= 8'b00000000 ;
			15'h0000190D : data <= 8'b00000000 ;
			15'h0000190E : data <= 8'b00000000 ;
			15'h0000190F : data <= 8'b00000000 ;
			15'h00001910 : data <= 8'b00000000 ;
			15'h00001911 : data <= 8'b00000000 ;
			15'h00001912 : data <= 8'b00000000 ;
			15'h00001913 : data <= 8'b00000000 ;
			15'h00001914 : data <= 8'b00000000 ;
			15'h00001915 : data <= 8'b00000000 ;
			15'h00001916 : data <= 8'b00000000 ;
			15'h00001917 : data <= 8'b00000000 ;
			15'h00001918 : data <= 8'b00000000 ;
			15'h00001919 : data <= 8'b00000000 ;
			15'h0000191A : data <= 8'b00000000 ;
			15'h0000191B : data <= 8'b00000000 ;
			15'h0000191C : data <= 8'b00000000 ;
			15'h0000191D : data <= 8'b00000000 ;
			15'h0000191E : data <= 8'b00000000 ;
			15'h0000191F : data <= 8'b00000000 ;
			15'h00001920 : data <= 8'b00000000 ;
			15'h00001921 : data <= 8'b00000000 ;
			15'h00001922 : data <= 8'b00000000 ;
			15'h00001923 : data <= 8'b00000000 ;
			15'h00001924 : data <= 8'b00000000 ;
			15'h00001925 : data <= 8'b00000000 ;
			15'h00001926 : data <= 8'b00000000 ;
			15'h00001927 : data <= 8'b00000000 ;
			15'h00001928 : data <= 8'b00000000 ;
			15'h00001929 : data <= 8'b00000000 ;
			15'h0000192A : data <= 8'b00000000 ;
			15'h0000192B : data <= 8'b00000000 ;
			15'h0000192C : data <= 8'b00000000 ;
			15'h0000192D : data <= 8'b00000000 ;
			15'h0000192E : data <= 8'b00000000 ;
			15'h0000192F : data <= 8'b00000000 ;
			15'h00001930 : data <= 8'b00000000 ;
			15'h00001931 : data <= 8'b00000000 ;
			15'h00001932 : data <= 8'b00000000 ;
			15'h00001933 : data <= 8'b00000000 ;
			15'h00001934 : data <= 8'b00000000 ;
			15'h00001935 : data <= 8'b00000000 ;
			15'h00001936 : data <= 8'b00000000 ;
			15'h00001937 : data <= 8'b00000000 ;
			15'h00001938 : data <= 8'b00000000 ;
			15'h00001939 : data <= 8'b00000000 ;
			15'h0000193A : data <= 8'b00000000 ;
			15'h0000193B : data <= 8'b00000000 ;
			15'h0000193C : data <= 8'b00000000 ;
			15'h0000193D : data <= 8'b00000000 ;
			15'h0000193E : data <= 8'b00000000 ;
			15'h0000193F : data <= 8'b00000000 ;
			15'h00001940 : data <= 8'b00000000 ;
			15'h00001941 : data <= 8'b00000000 ;
			15'h00001942 : data <= 8'b00000000 ;
			15'h00001943 : data <= 8'b00000000 ;
			15'h00001944 : data <= 8'b00000000 ;
			15'h00001945 : data <= 8'b00000000 ;
			15'h00001946 : data <= 8'b00000000 ;
			15'h00001947 : data <= 8'b00000000 ;
			15'h00001948 : data <= 8'b00000000 ;
			15'h00001949 : data <= 8'b00000000 ;
			15'h0000194A : data <= 8'b00000000 ;
			15'h0000194B : data <= 8'b00000000 ;
			15'h0000194C : data <= 8'b00000000 ;
			15'h0000194D : data <= 8'b00000000 ;
			15'h0000194E : data <= 8'b00000000 ;
			15'h0000194F : data <= 8'b00000000 ;
			15'h00001950 : data <= 8'b00000000 ;
			15'h00001951 : data <= 8'b00000000 ;
			15'h00001952 : data <= 8'b00000000 ;
			15'h00001953 : data <= 8'b00000000 ;
			15'h00001954 : data <= 8'b00000000 ;
			15'h00001955 : data <= 8'b00000000 ;
			15'h00001956 : data <= 8'b00000000 ;
			15'h00001957 : data <= 8'b00000000 ;
			15'h00001958 : data <= 8'b00000000 ;
			15'h00001959 : data <= 8'b00000000 ;
			15'h0000195A : data <= 8'b00000000 ;
			15'h0000195B : data <= 8'b00000000 ;
			15'h0000195C : data <= 8'b00000000 ;
			15'h0000195D : data <= 8'b00000000 ;
			15'h0000195E : data <= 8'b00000000 ;
			15'h0000195F : data <= 8'b00000000 ;
			15'h00001960 : data <= 8'b00000000 ;
			15'h00001961 : data <= 8'b00000000 ;
			15'h00001962 : data <= 8'b00000000 ;
			15'h00001963 : data <= 8'b00000000 ;
			15'h00001964 : data <= 8'b00000000 ;
			15'h00001965 : data <= 8'b00000000 ;
			15'h00001966 : data <= 8'b00000000 ;
			15'h00001967 : data <= 8'b00000000 ;
			15'h00001968 : data <= 8'b00000000 ;
			15'h00001969 : data <= 8'b00000000 ;
			15'h0000196A : data <= 8'b00000000 ;
			15'h0000196B : data <= 8'b00000000 ;
			15'h0000196C : data <= 8'b00000000 ;
			15'h0000196D : data <= 8'b00000000 ;
			15'h0000196E : data <= 8'b00000000 ;
			15'h0000196F : data <= 8'b00000000 ;
			15'h00001970 : data <= 8'b00000000 ;
			15'h00001971 : data <= 8'b00000000 ;
			15'h00001972 : data <= 8'b00000000 ;
			15'h00001973 : data <= 8'b00000000 ;
			15'h00001974 : data <= 8'b00000000 ;
			15'h00001975 : data <= 8'b00000000 ;
			15'h00001976 : data <= 8'b00000000 ;
			15'h00001977 : data <= 8'b00000000 ;
			15'h00001978 : data <= 8'b00000000 ;
			15'h00001979 : data <= 8'b00000000 ;
			15'h0000197A : data <= 8'b00000000 ;
			15'h0000197B : data <= 8'b00000000 ;
			15'h0000197C : data <= 8'b00000000 ;
			15'h0000197D : data <= 8'b00000000 ;
			15'h0000197E : data <= 8'b00000000 ;
			15'h0000197F : data <= 8'b00000000 ;
			15'h00001980 : data <= 8'b00000000 ;
			15'h00001981 : data <= 8'b00000000 ;
			15'h00001982 : data <= 8'b00000000 ;
			15'h00001983 : data <= 8'b00000000 ;
			15'h00001984 : data <= 8'b00000000 ;
			15'h00001985 : data <= 8'b00000000 ;
			15'h00001986 : data <= 8'b00000000 ;
			15'h00001987 : data <= 8'b00000000 ;
			15'h00001988 : data <= 8'b00000000 ;
			15'h00001989 : data <= 8'b00000000 ;
			15'h0000198A : data <= 8'b00000000 ;
			15'h0000198B : data <= 8'b00000000 ;
			15'h0000198C : data <= 8'b00000000 ;
			15'h0000198D : data <= 8'b00000000 ;
			15'h0000198E : data <= 8'b00000000 ;
			15'h0000198F : data <= 8'b00000000 ;
			15'h00001990 : data <= 8'b00000000 ;
			15'h00001991 : data <= 8'b00000000 ;
			15'h00001992 : data <= 8'b00000000 ;
			15'h00001993 : data <= 8'b00000000 ;
			15'h00001994 : data <= 8'b00000000 ;
			15'h00001995 : data <= 8'b00000000 ;
			15'h00001996 : data <= 8'b00000000 ;
			15'h00001997 : data <= 8'b00000000 ;
			15'h00001998 : data <= 8'b00000000 ;
			15'h00001999 : data <= 8'b00000000 ;
			15'h0000199A : data <= 8'b00000000 ;
			15'h0000199B : data <= 8'b00000000 ;
			15'h0000199C : data <= 8'b00000000 ;
			15'h0000199D : data <= 8'b00000000 ;
			15'h0000199E : data <= 8'b00000000 ;
			15'h0000199F : data <= 8'b00000000 ;
			15'h000019A0 : data <= 8'b00000000 ;
			15'h000019A1 : data <= 8'b00000000 ;
			15'h000019A2 : data <= 8'b00000000 ;
			15'h000019A3 : data <= 8'b00000000 ;
			15'h000019A4 : data <= 8'b00000000 ;
			15'h000019A5 : data <= 8'b00000000 ;
			15'h000019A6 : data <= 8'b00000000 ;
			15'h000019A7 : data <= 8'b00000000 ;
			15'h000019A8 : data <= 8'b00000000 ;
			15'h000019A9 : data <= 8'b00000000 ;
			15'h000019AA : data <= 8'b00000000 ;
			15'h000019AB : data <= 8'b00000000 ;
			15'h000019AC : data <= 8'b00000000 ;
			15'h000019AD : data <= 8'b00000000 ;
			15'h000019AE : data <= 8'b00000000 ;
			15'h000019AF : data <= 8'b00000000 ;
			15'h000019B0 : data <= 8'b00000000 ;
			15'h000019B1 : data <= 8'b00000000 ;
			15'h000019B2 : data <= 8'b00000000 ;
			15'h000019B3 : data <= 8'b00000000 ;
			15'h000019B4 : data <= 8'b00000000 ;
			15'h000019B5 : data <= 8'b00000000 ;
			15'h000019B6 : data <= 8'b00000000 ;
			15'h000019B7 : data <= 8'b00000000 ;
			15'h000019B8 : data <= 8'b00000000 ;
			15'h000019B9 : data <= 8'b00000000 ;
			15'h000019BA : data <= 8'b00000000 ;
			15'h000019BB : data <= 8'b00000000 ;
			15'h000019BC : data <= 8'b00000000 ;
			15'h000019BD : data <= 8'b00000000 ;
			15'h000019BE : data <= 8'b00000000 ;
			15'h000019BF : data <= 8'b00000000 ;
			15'h000019C0 : data <= 8'b00000000 ;
			15'h000019C1 : data <= 8'b00000000 ;
			15'h000019C2 : data <= 8'b00000000 ;
			15'h000019C3 : data <= 8'b00000000 ;
			15'h000019C4 : data <= 8'b00000000 ;
			15'h000019C5 : data <= 8'b00000000 ;
			15'h000019C6 : data <= 8'b00000000 ;
			15'h000019C7 : data <= 8'b00000000 ;
			15'h000019C8 : data <= 8'b00000000 ;
			15'h000019C9 : data <= 8'b00000000 ;
			15'h000019CA : data <= 8'b00000000 ;
			15'h000019CB : data <= 8'b00000000 ;
			15'h000019CC : data <= 8'b00000000 ;
			15'h000019CD : data <= 8'b00000000 ;
			15'h000019CE : data <= 8'b00000000 ;
			15'h000019CF : data <= 8'b00000000 ;
			15'h000019D0 : data <= 8'b00000000 ;
			15'h000019D1 : data <= 8'b00000000 ;
			15'h000019D2 : data <= 8'b00000000 ;
			15'h000019D3 : data <= 8'b00000000 ;
			15'h000019D4 : data <= 8'b00000000 ;
			15'h000019D5 : data <= 8'b00000000 ;
			15'h000019D6 : data <= 8'b00000000 ;
			15'h000019D7 : data <= 8'b00000000 ;
			15'h000019D8 : data <= 8'b00000000 ;
			15'h000019D9 : data <= 8'b00000000 ;
			15'h000019DA : data <= 8'b00000000 ;
			15'h000019DB : data <= 8'b00000000 ;
			15'h000019DC : data <= 8'b00000000 ;
			15'h000019DD : data <= 8'b00000000 ;
			15'h000019DE : data <= 8'b00000000 ;
			15'h000019DF : data <= 8'b00000000 ;
			15'h000019E0 : data <= 8'b00000000 ;
			15'h000019E1 : data <= 8'b00000000 ;
			15'h000019E2 : data <= 8'b00000000 ;
			15'h000019E3 : data <= 8'b00000000 ;
			15'h000019E4 : data <= 8'b00000000 ;
			15'h000019E5 : data <= 8'b00000000 ;
			15'h000019E6 : data <= 8'b00000000 ;
			15'h000019E7 : data <= 8'b00000000 ;
			15'h000019E8 : data <= 8'b00000000 ;
			15'h000019E9 : data <= 8'b00000000 ;
			15'h000019EA : data <= 8'b00000000 ;
			15'h000019EB : data <= 8'b00000000 ;
			15'h000019EC : data <= 8'b00000000 ;
			15'h000019ED : data <= 8'b00000000 ;
			15'h000019EE : data <= 8'b00000000 ;
			15'h000019EF : data <= 8'b00000000 ;
			15'h000019F0 : data <= 8'b00000000 ;
			15'h000019F1 : data <= 8'b00000000 ;
			15'h000019F2 : data <= 8'b00000000 ;
			15'h000019F3 : data <= 8'b00000000 ;
			15'h000019F4 : data <= 8'b00000000 ;
			15'h000019F5 : data <= 8'b00000000 ;
			15'h000019F6 : data <= 8'b00000000 ;
			15'h000019F7 : data <= 8'b00000000 ;
			15'h000019F8 : data <= 8'b00000000 ;
			15'h000019F9 : data <= 8'b00000000 ;
			15'h000019FA : data <= 8'b00000000 ;
			15'h000019FB : data <= 8'b00000000 ;
			15'h000019FC : data <= 8'b00000000 ;
			15'h000019FD : data <= 8'b00000000 ;
			15'h000019FE : data <= 8'b00000000 ;
			15'h000019FF : data <= 8'b00000000 ;
			15'h00001A00 : data <= 8'b00000000 ;
			15'h00001A01 : data <= 8'b00000000 ;
			15'h00001A02 : data <= 8'b00000000 ;
			15'h00001A03 : data <= 8'b00000000 ;
			15'h00001A04 : data <= 8'b00000000 ;
			15'h00001A05 : data <= 8'b00000000 ;
			15'h00001A06 : data <= 8'b00000000 ;
			15'h00001A07 : data <= 8'b00000000 ;
			15'h00001A08 : data <= 8'b00000000 ;
			15'h00001A09 : data <= 8'b00000000 ;
			15'h00001A0A : data <= 8'b00000000 ;
			15'h00001A0B : data <= 8'b00000000 ;
			15'h00001A0C : data <= 8'b00000000 ;
			15'h00001A0D : data <= 8'b00000000 ;
			15'h00001A0E : data <= 8'b00000000 ;
			15'h00001A0F : data <= 8'b00000000 ;
			15'h00001A10 : data <= 8'b00000000 ;
			15'h00001A11 : data <= 8'b00000000 ;
			15'h00001A12 : data <= 8'b00000000 ;
			15'h00001A13 : data <= 8'b00000000 ;
			15'h00001A14 : data <= 8'b00000000 ;
			15'h00001A15 : data <= 8'b00000000 ;
			15'h00001A16 : data <= 8'b00000000 ;
			15'h00001A17 : data <= 8'b00000000 ;
			15'h00001A18 : data <= 8'b00000000 ;
			15'h00001A19 : data <= 8'b00000000 ;
			15'h00001A1A : data <= 8'b00000000 ;
			15'h00001A1B : data <= 8'b00000000 ;
			15'h00001A1C : data <= 8'b00000000 ;
			15'h00001A1D : data <= 8'b00000000 ;
			15'h00001A1E : data <= 8'b00000000 ;
			15'h00001A1F : data <= 8'b00000000 ;
			15'h00001A20 : data <= 8'b00000000 ;
			15'h00001A21 : data <= 8'b00000000 ;
			15'h00001A22 : data <= 8'b00000000 ;
			15'h00001A23 : data <= 8'b00000000 ;
			15'h00001A24 : data <= 8'b00000000 ;
			15'h00001A25 : data <= 8'b00000000 ;
			15'h00001A26 : data <= 8'b00000000 ;
			15'h00001A27 : data <= 8'b00000000 ;
			15'h00001A28 : data <= 8'b00000000 ;
			15'h00001A29 : data <= 8'b00000000 ;
			15'h00001A2A : data <= 8'b00000000 ;
			15'h00001A2B : data <= 8'b00000000 ;
			15'h00001A2C : data <= 8'b00000000 ;
			15'h00001A2D : data <= 8'b00000000 ;
			15'h00001A2E : data <= 8'b00000000 ;
			15'h00001A2F : data <= 8'b00000000 ;
			15'h00001A30 : data <= 8'b00000000 ;
			15'h00001A31 : data <= 8'b00000000 ;
			15'h00001A32 : data <= 8'b00000000 ;
			15'h00001A33 : data <= 8'b00000000 ;
			15'h00001A34 : data <= 8'b00000000 ;
			15'h00001A35 : data <= 8'b00000000 ;
			15'h00001A36 : data <= 8'b00000000 ;
			15'h00001A37 : data <= 8'b00000000 ;
			15'h00001A38 : data <= 8'b00000000 ;
			15'h00001A39 : data <= 8'b00000000 ;
			15'h00001A3A : data <= 8'b00000000 ;
			15'h00001A3B : data <= 8'b00000000 ;
			15'h00001A3C : data <= 8'b00000000 ;
			15'h00001A3D : data <= 8'b00000000 ;
			15'h00001A3E : data <= 8'b00000000 ;
			15'h00001A3F : data <= 8'b00000000 ;
			15'h00001A40 : data <= 8'b00000000 ;
			15'h00001A41 : data <= 8'b00000000 ;
			15'h00001A42 : data <= 8'b00000000 ;
			15'h00001A43 : data <= 8'b00000000 ;
			15'h00001A44 : data <= 8'b00000000 ;
			15'h00001A45 : data <= 8'b00000000 ;
			15'h00001A46 : data <= 8'b00000000 ;
			15'h00001A47 : data <= 8'b00000000 ;
			15'h00001A48 : data <= 8'b00000000 ;
			15'h00001A49 : data <= 8'b00000000 ;
			15'h00001A4A : data <= 8'b00000000 ;
			15'h00001A4B : data <= 8'b00000000 ;
			15'h00001A4C : data <= 8'b00000000 ;
			15'h00001A4D : data <= 8'b00000000 ;
			15'h00001A4E : data <= 8'b00000000 ;
			15'h00001A4F : data <= 8'b00000000 ;
			15'h00001A50 : data <= 8'b00000000 ;
			15'h00001A51 : data <= 8'b00000000 ;
			15'h00001A52 : data <= 8'b00000000 ;
			15'h00001A53 : data <= 8'b00000000 ;
			15'h00001A54 : data <= 8'b00000000 ;
			15'h00001A55 : data <= 8'b00000000 ;
			15'h00001A56 : data <= 8'b00000000 ;
			15'h00001A57 : data <= 8'b00000000 ;
			15'h00001A58 : data <= 8'b00000000 ;
			15'h00001A59 : data <= 8'b00000000 ;
			15'h00001A5A : data <= 8'b00000000 ;
			15'h00001A5B : data <= 8'b00000000 ;
			15'h00001A5C : data <= 8'b00000000 ;
			15'h00001A5D : data <= 8'b00000000 ;
			15'h00001A5E : data <= 8'b00000000 ;
			15'h00001A5F : data <= 8'b00000000 ;
			15'h00001A60 : data <= 8'b00000000 ;
			15'h00001A61 : data <= 8'b00000000 ;
			15'h00001A62 : data <= 8'b00000000 ;
			15'h00001A63 : data <= 8'b00000000 ;
			15'h00001A64 : data <= 8'b00000000 ;
			15'h00001A65 : data <= 8'b00000000 ;
			15'h00001A66 : data <= 8'b00000000 ;
			15'h00001A67 : data <= 8'b00000000 ;
			15'h00001A68 : data <= 8'b00000000 ;
			15'h00001A69 : data <= 8'b00000000 ;
			15'h00001A6A : data <= 8'b00000000 ;
			15'h00001A6B : data <= 8'b00000000 ;
			15'h00001A6C : data <= 8'b00000000 ;
			15'h00001A6D : data <= 8'b00000000 ;
			15'h00001A6E : data <= 8'b00000000 ;
			15'h00001A6F : data <= 8'b00000000 ;
			15'h00001A70 : data <= 8'b00000000 ;
			15'h00001A71 : data <= 8'b00000000 ;
			15'h00001A72 : data <= 8'b00000000 ;
			15'h00001A73 : data <= 8'b00000000 ;
			15'h00001A74 : data <= 8'b00000000 ;
			15'h00001A75 : data <= 8'b00000000 ;
			15'h00001A76 : data <= 8'b00000000 ;
			15'h00001A77 : data <= 8'b00000000 ;
			15'h00001A78 : data <= 8'b00000000 ;
			15'h00001A79 : data <= 8'b00000000 ;
			15'h00001A7A : data <= 8'b00000000 ;
			15'h00001A7B : data <= 8'b00000000 ;
			15'h00001A7C : data <= 8'b00000000 ;
			15'h00001A7D : data <= 8'b00000000 ;
			15'h00001A7E : data <= 8'b00000000 ;
			15'h00001A7F : data <= 8'b00000000 ;
			15'h00001A80 : data <= 8'b00000000 ;
			15'h00001A81 : data <= 8'b00000000 ;
			15'h00001A82 : data <= 8'b00000000 ;
			15'h00001A83 : data <= 8'b00000000 ;
			15'h00001A84 : data <= 8'b00000000 ;
			15'h00001A85 : data <= 8'b00000000 ;
			15'h00001A86 : data <= 8'b00000000 ;
			15'h00001A87 : data <= 8'b00000000 ;
			15'h00001A88 : data <= 8'b00000000 ;
			15'h00001A89 : data <= 8'b00000000 ;
			15'h00001A8A : data <= 8'b00000000 ;
			15'h00001A8B : data <= 8'b00000000 ;
			15'h00001A8C : data <= 8'b00000000 ;
			15'h00001A8D : data <= 8'b00000000 ;
			15'h00001A8E : data <= 8'b00000000 ;
			15'h00001A8F : data <= 8'b00000000 ;
			15'h00001A90 : data <= 8'b00000000 ;
			15'h00001A91 : data <= 8'b00000000 ;
			15'h00001A92 : data <= 8'b00000000 ;
			15'h00001A93 : data <= 8'b00000000 ;
			15'h00001A94 : data <= 8'b00000000 ;
			15'h00001A95 : data <= 8'b00000000 ;
			15'h00001A96 : data <= 8'b00000000 ;
			15'h00001A97 : data <= 8'b00000000 ;
			15'h00001A98 : data <= 8'b00000000 ;
			15'h00001A99 : data <= 8'b00000000 ;
			15'h00001A9A : data <= 8'b00000000 ;
			15'h00001A9B : data <= 8'b00000000 ;
			15'h00001A9C : data <= 8'b00000000 ;
			15'h00001A9D : data <= 8'b00000000 ;
			15'h00001A9E : data <= 8'b00000000 ;
			15'h00001A9F : data <= 8'b00000000 ;
			15'h00001AA0 : data <= 8'b00000000 ;
			15'h00001AA1 : data <= 8'b00000000 ;
			15'h00001AA2 : data <= 8'b00000000 ;
			15'h00001AA3 : data <= 8'b00000000 ;
			15'h00001AA4 : data <= 8'b00000000 ;
			15'h00001AA5 : data <= 8'b00000000 ;
			15'h00001AA6 : data <= 8'b00000000 ;
			15'h00001AA7 : data <= 8'b00000000 ;
			15'h00001AA8 : data <= 8'b00000000 ;
			15'h00001AA9 : data <= 8'b00000000 ;
			15'h00001AAA : data <= 8'b00000000 ;
			15'h00001AAB : data <= 8'b00000000 ;
			15'h00001AAC : data <= 8'b00000000 ;
			15'h00001AAD : data <= 8'b00000000 ;
			15'h00001AAE : data <= 8'b00000000 ;
			15'h00001AAF : data <= 8'b00000000 ;
			15'h00001AB0 : data <= 8'b00000000 ;
			15'h00001AB1 : data <= 8'b00000000 ;
			15'h00001AB2 : data <= 8'b00000000 ;
			15'h00001AB3 : data <= 8'b00000000 ;
			15'h00001AB4 : data <= 8'b00000000 ;
			15'h00001AB5 : data <= 8'b00000000 ;
			15'h00001AB6 : data <= 8'b00000000 ;
			15'h00001AB7 : data <= 8'b00000000 ;
			15'h00001AB8 : data <= 8'b00000000 ;
			15'h00001AB9 : data <= 8'b00000000 ;
			15'h00001ABA : data <= 8'b00000000 ;
			15'h00001ABB : data <= 8'b00000000 ;
			15'h00001ABC : data <= 8'b00000000 ;
			15'h00001ABD : data <= 8'b00000000 ;
			15'h00001ABE : data <= 8'b00000000 ;
			15'h00001ABF : data <= 8'b00000000 ;
			15'h00001AC0 : data <= 8'b00000000 ;
			15'h00001AC1 : data <= 8'b00000000 ;
			15'h00001AC2 : data <= 8'b00000000 ;
			15'h00001AC3 : data <= 8'b00000000 ;
			15'h00001AC4 : data <= 8'b00000000 ;
			15'h00001AC5 : data <= 8'b00000000 ;
			15'h00001AC6 : data <= 8'b00000000 ;
			15'h00001AC7 : data <= 8'b00000000 ;
			15'h00001AC8 : data <= 8'b00000000 ;
			15'h00001AC9 : data <= 8'b00000000 ;
			15'h00001ACA : data <= 8'b00000000 ;
			15'h00001ACB : data <= 8'b00000000 ;
			15'h00001ACC : data <= 8'b00000000 ;
			15'h00001ACD : data <= 8'b00000000 ;
			15'h00001ACE : data <= 8'b00000000 ;
			15'h00001ACF : data <= 8'b00000000 ;
			15'h00001AD0 : data <= 8'b00000000 ;
			15'h00001AD1 : data <= 8'b00000000 ;
			15'h00001AD2 : data <= 8'b00000000 ;
			15'h00001AD3 : data <= 8'b00000000 ;
			15'h00001AD4 : data <= 8'b00000000 ;
			15'h00001AD5 : data <= 8'b00000000 ;
			15'h00001AD6 : data <= 8'b00000000 ;
			15'h00001AD7 : data <= 8'b00000000 ;
			15'h00001AD8 : data <= 8'b00000000 ;
			15'h00001AD9 : data <= 8'b00000000 ;
			15'h00001ADA : data <= 8'b00000000 ;
			15'h00001ADB : data <= 8'b00000000 ;
			15'h00001ADC : data <= 8'b00000000 ;
			15'h00001ADD : data <= 8'b00000000 ;
			15'h00001ADE : data <= 8'b00000000 ;
			15'h00001ADF : data <= 8'b00000000 ;
			15'h00001AE0 : data <= 8'b00000000 ;
			15'h00001AE1 : data <= 8'b00000000 ;
			15'h00001AE2 : data <= 8'b00000000 ;
			15'h00001AE3 : data <= 8'b00000000 ;
			15'h00001AE4 : data <= 8'b00000000 ;
			15'h00001AE5 : data <= 8'b00000000 ;
			15'h00001AE6 : data <= 8'b00000000 ;
			15'h00001AE7 : data <= 8'b00000000 ;
			15'h00001AE8 : data <= 8'b00000000 ;
			15'h00001AE9 : data <= 8'b00000000 ;
			15'h00001AEA : data <= 8'b00000000 ;
			15'h00001AEB : data <= 8'b00000000 ;
			15'h00001AEC : data <= 8'b00000000 ;
			15'h00001AED : data <= 8'b00000000 ;
			15'h00001AEE : data <= 8'b00000000 ;
			15'h00001AEF : data <= 8'b00000000 ;
			15'h00001AF0 : data <= 8'b00000000 ;
			15'h00001AF1 : data <= 8'b00000000 ;
			15'h00001AF2 : data <= 8'b00000000 ;
			15'h00001AF3 : data <= 8'b00000000 ;
			15'h00001AF4 : data <= 8'b00000000 ;
			15'h00001AF5 : data <= 8'b00000000 ;
			15'h00001AF6 : data <= 8'b00000000 ;
			15'h00001AF7 : data <= 8'b00000000 ;
			15'h00001AF8 : data <= 8'b00000000 ;
			15'h00001AF9 : data <= 8'b00000000 ;
			15'h00001AFA : data <= 8'b00000000 ;
			15'h00001AFB : data <= 8'b00000000 ;
			15'h00001AFC : data <= 8'b00000000 ;
			15'h00001AFD : data <= 8'b00000000 ;
			15'h00001AFE : data <= 8'b00000000 ;
			15'h00001AFF : data <= 8'b00000000 ;
			15'h00001B00 : data <= 8'b00000000 ;
			15'h00001B01 : data <= 8'b00000000 ;
			15'h00001B02 : data <= 8'b00000000 ;
			15'h00001B03 : data <= 8'b00000000 ;
			15'h00001B04 : data <= 8'b00000000 ;
			15'h00001B05 : data <= 8'b00000000 ;
			15'h00001B06 : data <= 8'b00000000 ;
			15'h00001B07 : data <= 8'b00000000 ;
			15'h00001B08 : data <= 8'b00000000 ;
			15'h00001B09 : data <= 8'b00000000 ;
			15'h00001B0A : data <= 8'b00000000 ;
			15'h00001B0B : data <= 8'b00000000 ;
			15'h00001B0C : data <= 8'b00000000 ;
			15'h00001B0D : data <= 8'b00000000 ;
			15'h00001B0E : data <= 8'b00000000 ;
			15'h00001B0F : data <= 8'b00000000 ;
			15'h00001B10 : data <= 8'b00000000 ;
			15'h00001B11 : data <= 8'b00000000 ;
			15'h00001B12 : data <= 8'b00000000 ;
			15'h00001B13 : data <= 8'b00000000 ;
			15'h00001B14 : data <= 8'b00000000 ;
			15'h00001B15 : data <= 8'b00000000 ;
			15'h00001B16 : data <= 8'b00000000 ;
			15'h00001B17 : data <= 8'b00000000 ;
			15'h00001B18 : data <= 8'b00000000 ;
			15'h00001B19 : data <= 8'b00000000 ;
			15'h00001B1A : data <= 8'b00000000 ;
			15'h00001B1B : data <= 8'b00000000 ;
			15'h00001B1C : data <= 8'b00000000 ;
			15'h00001B1D : data <= 8'b00000000 ;
			15'h00001B1E : data <= 8'b00000000 ;
			15'h00001B1F : data <= 8'b00000000 ;
			15'h00001B20 : data <= 8'b00000000 ;
			15'h00001B21 : data <= 8'b00000000 ;
			15'h00001B22 : data <= 8'b00000000 ;
			15'h00001B23 : data <= 8'b00000000 ;
			15'h00001B24 : data <= 8'b00000000 ;
			15'h00001B25 : data <= 8'b00000000 ;
			15'h00001B26 : data <= 8'b00000000 ;
			15'h00001B27 : data <= 8'b00000000 ;
			15'h00001B28 : data <= 8'b00000000 ;
			15'h00001B29 : data <= 8'b00000000 ;
			15'h00001B2A : data <= 8'b00000000 ;
			15'h00001B2B : data <= 8'b00000000 ;
			15'h00001B2C : data <= 8'b00000000 ;
			15'h00001B2D : data <= 8'b00000000 ;
			15'h00001B2E : data <= 8'b00000000 ;
			15'h00001B2F : data <= 8'b00000000 ;
			15'h00001B30 : data <= 8'b00000000 ;
			15'h00001B31 : data <= 8'b00000000 ;
			15'h00001B32 : data <= 8'b00000000 ;
			15'h00001B33 : data <= 8'b00000000 ;
			15'h00001B34 : data <= 8'b00000000 ;
			15'h00001B35 : data <= 8'b00000000 ;
			15'h00001B36 : data <= 8'b00000000 ;
			15'h00001B37 : data <= 8'b00000000 ;
			15'h00001B38 : data <= 8'b00000000 ;
			15'h00001B39 : data <= 8'b00000000 ;
			15'h00001B3A : data <= 8'b00000000 ;
			15'h00001B3B : data <= 8'b00000000 ;
			15'h00001B3C : data <= 8'b00000000 ;
			15'h00001B3D : data <= 8'b00000000 ;
			15'h00001B3E : data <= 8'b00000000 ;
			15'h00001B3F : data <= 8'b00000000 ;
			15'h00001B40 : data <= 8'b00000000 ;
			15'h00001B41 : data <= 8'b00000000 ;
			15'h00001B42 : data <= 8'b00000000 ;
			15'h00001B43 : data <= 8'b00000000 ;
			15'h00001B44 : data <= 8'b00000000 ;
			15'h00001B45 : data <= 8'b00000000 ;
			15'h00001B46 : data <= 8'b00000000 ;
			15'h00001B47 : data <= 8'b00000000 ;
			15'h00001B48 : data <= 8'b00000000 ;
			15'h00001B49 : data <= 8'b00000000 ;
			15'h00001B4A : data <= 8'b00000000 ;
			15'h00001B4B : data <= 8'b00000000 ;
			15'h00001B4C : data <= 8'b00000000 ;
			15'h00001B4D : data <= 8'b00000000 ;
			15'h00001B4E : data <= 8'b00000000 ;
			15'h00001B4F : data <= 8'b00000000 ;
			15'h00001B50 : data <= 8'b00000000 ;
			15'h00001B51 : data <= 8'b00000000 ;
			15'h00001B52 : data <= 8'b00000000 ;
			15'h00001B53 : data <= 8'b00000000 ;
			15'h00001B54 : data <= 8'b00000000 ;
			15'h00001B55 : data <= 8'b00000000 ;
			15'h00001B56 : data <= 8'b00000000 ;
			15'h00001B57 : data <= 8'b00000000 ;
			15'h00001B58 : data <= 8'b00000000 ;
			15'h00001B59 : data <= 8'b00000000 ;
			15'h00001B5A : data <= 8'b00000000 ;
			15'h00001B5B : data <= 8'b00000000 ;
			15'h00001B5C : data <= 8'b00000000 ;
			15'h00001B5D : data <= 8'b00000000 ;
			15'h00001B5E : data <= 8'b00000000 ;
			15'h00001B5F : data <= 8'b00000000 ;
			15'h00001B60 : data <= 8'b00000000 ;
			15'h00001B61 : data <= 8'b00000000 ;
			15'h00001B62 : data <= 8'b00000000 ;
			15'h00001B63 : data <= 8'b00000000 ;
			15'h00001B64 : data <= 8'b00000000 ;
			15'h00001B65 : data <= 8'b00000000 ;
			15'h00001B66 : data <= 8'b00000000 ;
			15'h00001B67 : data <= 8'b00000000 ;
			15'h00001B68 : data <= 8'b00000000 ;
			15'h00001B69 : data <= 8'b00000000 ;
			15'h00001B6A : data <= 8'b00000000 ;
			15'h00001B6B : data <= 8'b00000000 ;
			15'h00001B6C : data <= 8'b00000000 ;
			15'h00001B6D : data <= 8'b00000000 ;
			15'h00001B6E : data <= 8'b00000000 ;
			15'h00001B6F : data <= 8'b00000000 ;
			15'h00001B70 : data <= 8'b00000000 ;
			15'h00001B71 : data <= 8'b00000000 ;
			15'h00001B72 : data <= 8'b00000000 ;
			15'h00001B73 : data <= 8'b00000000 ;
			15'h00001B74 : data <= 8'b00000000 ;
			15'h00001B75 : data <= 8'b00000000 ;
			15'h00001B76 : data <= 8'b00000000 ;
			15'h00001B77 : data <= 8'b00000000 ;
			15'h00001B78 : data <= 8'b00000000 ;
			15'h00001B79 : data <= 8'b00000000 ;
			15'h00001B7A : data <= 8'b00000000 ;
			15'h00001B7B : data <= 8'b00000000 ;
			15'h00001B7C : data <= 8'b00000000 ;
			15'h00001B7D : data <= 8'b00000000 ;
			15'h00001B7E : data <= 8'b00000000 ;
			15'h00001B7F : data <= 8'b00000000 ;
			15'h00001B80 : data <= 8'b00000000 ;
			15'h00001B81 : data <= 8'b00000000 ;
			15'h00001B82 : data <= 8'b00000000 ;
			15'h00001B83 : data <= 8'b00000000 ;
			15'h00001B84 : data <= 8'b00000000 ;
			15'h00001B85 : data <= 8'b00000000 ;
			15'h00001B86 : data <= 8'b00000000 ;
			15'h00001B87 : data <= 8'b00000000 ;
			15'h00001B88 : data <= 8'b00000000 ;
			15'h00001B89 : data <= 8'b00000000 ;
			15'h00001B8A : data <= 8'b00000000 ;
			15'h00001B8B : data <= 8'b00000000 ;
			15'h00001B8C : data <= 8'b00000000 ;
			15'h00001B8D : data <= 8'b00000000 ;
			15'h00001B8E : data <= 8'b00000000 ;
			15'h00001B8F : data <= 8'b00000000 ;
			15'h00001B90 : data <= 8'b00000000 ;
			15'h00001B91 : data <= 8'b00000000 ;
			15'h00001B92 : data <= 8'b00000000 ;
			15'h00001B93 : data <= 8'b00000000 ;
			15'h00001B94 : data <= 8'b00000000 ;
			15'h00001B95 : data <= 8'b00000000 ;
			15'h00001B96 : data <= 8'b00000000 ;
			15'h00001B97 : data <= 8'b00000000 ;
			15'h00001B98 : data <= 8'b00000000 ;
			15'h00001B99 : data <= 8'b00000000 ;
			15'h00001B9A : data <= 8'b00000000 ;
			15'h00001B9B : data <= 8'b00000000 ;
			15'h00001B9C : data <= 8'b00000000 ;
			15'h00001B9D : data <= 8'b00000000 ;
			15'h00001B9E : data <= 8'b00000000 ;
			15'h00001B9F : data <= 8'b00000000 ;
			15'h00001BA0 : data <= 8'b00000000 ;
			15'h00001BA1 : data <= 8'b00000000 ;
			15'h00001BA2 : data <= 8'b00000000 ;
			15'h00001BA3 : data <= 8'b00000000 ;
			15'h00001BA4 : data <= 8'b00000000 ;
			15'h00001BA5 : data <= 8'b00000000 ;
			15'h00001BA6 : data <= 8'b00000000 ;
			15'h00001BA7 : data <= 8'b00000000 ;
			15'h00001BA8 : data <= 8'b00000000 ;
			15'h00001BA9 : data <= 8'b00000000 ;
			15'h00001BAA : data <= 8'b00000000 ;
			15'h00001BAB : data <= 8'b00000000 ;
			15'h00001BAC : data <= 8'b00000000 ;
			15'h00001BAD : data <= 8'b00000000 ;
			15'h00001BAE : data <= 8'b00000000 ;
			15'h00001BAF : data <= 8'b00000000 ;
			15'h00001BB0 : data <= 8'b00000000 ;
			15'h00001BB1 : data <= 8'b00000000 ;
			15'h00001BB2 : data <= 8'b00000000 ;
			15'h00001BB3 : data <= 8'b00000000 ;
			15'h00001BB4 : data <= 8'b00000000 ;
			15'h00001BB5 : data <= 8'b00000000 ;
			15'h00001BB6 : data <= 8'b00000000 ;
			15'h00001BB7 : data <= 8'b00000000 ;
			15'h00001BB8 : data <= 8'b00000000 ;
			15'h00001BB9 : data <= 8'b00000000 ;
			15'h00001BBA : data <= 8'b00000000 ;
			15'h00001BBB : data <= 8'b00000000 ;
			15'h00001BBC : data <= 8'b00000000 ;
			15'h00001BBD : data <= 8'b00000000 ;
			15'h00001BBE : data <= 8'b00000000 ;
			15'h00001BBF : data <= 8'b00000000 ;
			15'h00001BC0 : data <= 8'b00000000 ;
			15'h00001BC1 : data <= 8'b00000000 ;
			15'h00001BC2 : data <= 8'b00000000 ;
			15'h00001BC3 : data <= 8'b00000000 ;
			15'h00001BC4 : data <= 8'b00000000 ;
			15'h00001BC5 : data <= 8'b00000000 ;
			15'h00001BC6 : data <= 8'b00000000 ;
			15'h00001BC7 : data <= 8'b00000000 ;
			15'h00001BC8 : data <= 8'b00000000 ;
			15'h00001BC9 : data <= 8'b00000000 ;
			15'h00001BCA : data <= 8'b00000000 ;
			15'h00001BCB : data <= 8'b00000000 ;
			15'h00001BCC : data <= 8'b00000000 ;
			15'h00001BCD : data <= 8'b00000000 ;
			15'h00001BCE : data <= 8'b00000000 ;
			15'h00001BCF : data <= 8'b00000000 ;
			15'h00001BD0 : data <= 8'b00000000 ;
			15'h00001BD1 : data <= 8'b00000000 ;
			15'h00001BD2 : data <= 8'b00000000 ;
			15'h00001BD3 : data <= 8'b00000000 ;
			15'h00001BD4 : data <= 8'b00000000 ;
			15'h00001BD5 : data <= 8'b00000000 ;
			15'h00001BD6 : data <= 8'b00000000 ;
			15'h00001BD7 : data <= 8'b00000000 ;
			15'h00001BD8 : data <= 8'b00000000 ;
			15'h00001BD9 : data <= 8'b00000000 ;
			15'h00001BDA : data <= 8'b00000000 ;
			15'h00001BDB : data <= 8'b00000000 ;
			15'h00001BDC : data <= 8'b00000000 ;
			15'h00001BDD : data <= 8'b00000000 ;
			15'h00001BDE : data <= 8'b00000000 ;
			15'h00001BDF : data <= 8'b00000000 ;
			15'h00001BE0 : data <= 8'b00000000 ;
			15'h00001BE1 : data <= 8'b00000000 ;
			15'h00001BE2 : data <= 8'b00000000 ;
			15'h00001BE3 : data <= 8'b00000000 ;
			15'h00001BE4 : data <= 8'b00000000 ;
			15'h00001BE5 : data <= 8'b00000000 ;
			15'h00001BE6 : data <= 8'b00000000 ;
			15'h00001BE7 : data <= 8'b00000000 ;
			15'h00001BE8 : data <= 8'b00000000 ;
			15'h00001BE9 : data <= 8'b00000000 ;
			15'h00001BEA : data <= 8'b00000000 ;
			15'h00001BEB : data <= 8'b00000000 ;
			15'h00001BEC : data <= 8'b00000000 ;
			15'h00001BED : data <= 8'b00000000 ;
			15'h00001BEE : data <= 8'b00000000 ;
			15'h00001BEF : data <= 8'b00000000 ;
			15'h00001BF0 : data <= 8'b00000000 ;
			15'h00001BF1 : data <= 8'b00000000 ;
			15'h00001BF2 : data <= 8'b00000000 ;
			15'h00001BF3 : data <= 8'b00000000 ;
			15'h00001BF4 : data <= 8'b00000000 ;
			15'h00001BF5 : data <= 8'b00000000 ;
			15'h00001BF6 : data <= 8'b00000000 ;
			15'h00001BF7 : data <= 8'b00000000 ;
			15'h00001BF8 : data <= 8'b00000000 ;
			15'h00001BF9 : data <= 8'b00000000 ;
			15'h00001BFA : data <= 8'b00000000 ;
			15'h00001BFB : data <= 8'b00000000 ;
			15'h00001BFC : data <= 8'b00000000 ;
			15'h00001BFD : data <= 8'b00000000 ;
			15'h00001BFE : data <= 8'b00000000 ;
			15'h00001BFF : data <= 8'b00000000 ;
			15'h00001C00 : data <= 8'b00000000 ;
			15'h00001C01 : data <= 8'b00000000 ;
			15'h00001C02 : data <= 8'b00000000 ;
			15'h00001C03 : data <= 8'b00000000 ;
			15'h00001C04 : data <= 8'b00000000 ;
			15'h00001C05 : data <= 8'b00000000 ;
			15'h00001C06 : data <= 8'b00000000 ;
			15'h00001C07 : data <= 8'b00000000 ;
			15'h00001C08 : data <= 8'b00000000 ;
			15'h00001C09 : data <= 8'b00000000 ;
			15'h00001C0A : data <= 8'b00000000 ;
			15'h00001C0B : data <= 8'b00000000 ;
			15'h00001C0C : data <= 8'b00000000 ;
			15'h00001C0D : data <= 8'b00000000 ;
			15'h00001C0E : data <= 8'b00000000 ;
			15'h00001C0F : data <= 8'b00000000 ;
			15'h00001C10 : data <= 8'b00000000 ;
			15'h00001C11 : data <= 8'b00000000 ;
			15'h00001C12 : data <= 8'b00000000 ;
			15'h00001C13 : data <= 8'b00000000 ;
			15'h00001C14 : data <= 8'b00000000 ;
			15'h00001C15 : data <= 8'b00000000 ;
			15'h00001C16 : data <= 8'b00000000 ;
			15'h00001C17 : data <= 8'b00000000 ;
			15'h00001C18 : data <= 8'b00000000 ;
			15'h00001C19 : data <= 8'b00000000 ;
			15'h00001C1A : data <= 8'b00000000 ;
			15'h00001C1B : data <= 8'b00000000 ;
			15'h00001C1C : data <= 8'b00000000 ;
			15'h00001C1D : data <= 8'b00000000 ;
			15'h00001C1E : data <= 8'b00000000 ;
			15'h00001C1F : data <= 8'b00000000 ;
			15'h00001C20 : data <= 8'b00000000 ;
			15'h00001C21 : data <= 8'b00000000 ;
			15'h00001C22 : data <= 8'b00000000 ;
			15'h00001C23 : data <= 8'b00000000 ;
			15'h00001C24 : data <= 8'b00000000 ;
			15'h00001C25 : data <= 8'b00000000 ;
			15'h00001C26 : data <= 8'b00000000 ;
			15'h00001C27 : data <= 8'b00000000 ;
			15'h00001C28 : data <= 8'b00000000 ;
			15'h00001C29 : data <= 8'b00000000 ;
			15'h00001C2A : data <= 8'b00000000 ;
			15'h00001C2B : data <= 8'b00000000 ;
			15'h00001C2C : data <= 8'b00000000 ;
			15'h00001C2D : data <= 8'b00000000 ;
			15'h00001C2E : data <= 8'b00000000 ;
			15'h00001C2F : data <= 8'b00000000 ;
			15'h00001C30 : data <= 8'b00000000 ;
			15'h00001C31 : data <= 8'b00000000 ;
			15'h00001C32 : data <= 8'b00000000 ;
			15'h00001C33 : data <= 8'b00000000 ;
			15'h00001C34 : data <= 8'b00000000 ;
			15'h00001C35 : data <= 8'b00000000 ;
			15'h00001C36 : data <= 8'b00000000 ;
			15'h00001C37 : data <= 8'b00000000 ;
			15'h00001C38 : data <= 8'b00000000 ;
			15'h00001C39 : data <= 8'b00000000 ;
			15'h00001C3A : data <= 8'b00000000 ;
			15'h00001C3B : data <= 8'b00000000 ;
			15'h00001C3C : data <= 8'b00000000 ;
			15'h00001C3D : data <= 8'b00000000 ;
			15'h00001C3E : data <= 8'b00000000 ;
			15'h00001C3F : data <= 8'b00000000 ;
			15'h00001C40 : data <= 8'b00000000 ;
			15'h00001C41 : data <= 8'b00000000 ;
			15'h00001C42 : data <= 8'b00000000 ;
			15'h00001C43 : data <= 8'b00000000 ;
			15'h00001C44 : data <= 8'b00000000 ;
			15'h00001C45 : data <= 8'b00000000 ;
			15'h00001C46 : data <= 8'b00000000 ;
			15'h00001C47 : data <= 8'b00000000 ;
			15'h00001C48 : data <= 8'b00000000 ;
			15'h00001C49 : data <= 8'b00000000 ;
			15'h00001C4A : data <= 8'b00000000 ;
			15'h00001C4B : data <= 8'b00000000 ;
			15'h00001C4C : data <= 8'b00000000 ;
			15'h00001C4D : data <= 8'b00000000 ;
			15'h00001C4E : data <= 8'b00000000 ;
			15'h00001C4F : data <= 8'b00000000 ;
			15'h00001C50 : data <= 8'b00000000 ;
			15'h00001C51 : data <= 8'b00000000 ;
			15'h00001C52 : data <= 8'b00000000 ;
			15'h00001C53 : data <= 8'b00000000 ;
			15'h00001C54 : data <= 8'b00000000 ;
			15'h00001C55 : data <= 8'b00000000 ;
			15'h00001C56 : data <= 8'b00000000 ;
			15'h00001C57 : data <= 8'b00000000 ;
			15'h00001C58 : data <= 8'b00000000 ;
			15'h00001C59 : data <= 8'b00000000 ;
			15'h00001C5A : data <= 8'b00000000 ;
			15'h00001C5B : data <= 8'b00000000 ;
			15'h00001C5C : data <= 8'b00000000 ;
			15'h00001C5D : data <= 8'b00000000 ;
			15'h00001C5E : data <= 8'b00000000 ;
			15'h00001C5F : data <= 8'b00000000 ;
			15'h00001C60 : data <= 8'b00000000 ;
			15'h00001C61 : data <= 8'b00000000 ;
			15'h00001C62 : data <= 8'b00000000 ;
			15'h00001C63 : data <= 8'b00000000 ;
			15'h00001C64 : data <= 8'b00000000 ;
			15'h00001C65 : data <= 8'b00000000 ;
			15'h00001C66 : data <= 8'b00000000 ;
			15'h00001C67 : data <= 8'b00000000 ;
			15'h00001C68 : data <= 8'b00000000 ;
			15'h00001C69 : data <= 8'b00000000 ;
			15'h00001C6A : data <= 8'b00000000 ;
			15'h00001C6B : data <= 8'b00000000 ;
			15'h00001C6C : data <= 8'b00000000 ;
			15'h00001C6D : data <= 8'b00000000 ;
			15'h00001C6E : data <= 8'b00000000 ;
			15'h00001C6F : data <= 8'b00000000 ;
			15'h00001C70 : data <= 8'b00000000 ;
			15'h00001C71 : data <= 8'b00000000 ;
			15'h00001C72 : data <= 8'b00000000 ;
			15'h00001C73 : data <= 8'b00000000 ;
			15'h00001C74 : data <= 8'b00000000 ;
			15'h00001C75 : data <= 8'b00000000 ;
			15'h00001C76 : data <= 8'b00000000 ;
			15'h00001C77 : data <= 8'b00000000 ;
			15'h00001C78 : data <= 8'b00000000 ;
			15'h00001C79 : data <= 8'b00000000 ;
			15'h00001C7A : data <= 8'b00000000 ;
			15'h00001C7B : data <= 8'b00000000 ;
			15'h00001C7C : data <= 8'b00000000 ;
			15'h00001C7D : data <= 8'b00000000 ;
			15'h00001C7E : data <= 8'b00000000 ;
			15'h00001C7F : data <= 8'b00000000 ;
			15'h00001C80 : data <= 8'b00000000 ;
			15'h00001C81 : data <= 8'b00000000 ;
			15'h00001C82 : data <= 8'b00000000 ;
			15'h00001C83 : data <= 8'b00000000 ;
			15'h00001C84 : data <= 8'b00000000 ;
			15'h00001C85 : data <= 8'b00000000 ;
			15'h00001C86 : data <= 8'b00000000 ;
			15'h00001C87 : data <= 8'b00000000 ;
			15'h00001C88 : data <= 8'b00000000 ;
			15'h00001C89 : data <= 8'b00000000 ;
			15'h00001C8A : data <= 8'b00000000 ;
			15'h00001C8B : data <= 8'b00000000 ;
			15'h00001C8C : data <= 8'b00000000 ;
			15'h00001C8D : data <= 8'b00000000 ;
			15'h00001C8E : data <= 8'b00000000 ;
			15'h00001C8F : data <= 8'b00000000 ;
			15'h00001C90 : data <= 8'b00000000 ;
			15'h00001C91 : data <= 8'b00000000 ;
			15'h00001C92 : data <= 8'b00000000 ;
			15'h00001C93 : data <= 8'b00000000 ;
			15'h00001C94 : data <= 8'b00000000 ;
			15'h00001C95 : data <= 8'b00000000 ;
			15'h00001C96 : data <= 8'b00000000 ;
			15'h00001C97 : data <= 8'b00000000 ;
			15'h00001C98 : data <= 8'b00000000 ;
			15'h00001C99 : data <= 8'b00000000 ;
			15'h00001C9A : data <= 8'b00000000 ;
			15'h00001C9B : data <= 8'b00000000 ;
			15'h00001C9C : data <= 8'b00000000 ;
			15'h00001C9D : data <= 8'b00000000 ;
			15'h00001C9E : data <= 8'b00000000 ;
			15'h00001C9F : data <= 8'b00000000 ;
			15'h00001CA0 : data <= 8'b00000000 ;
			15'h00001CA1 : data <= 8'b00000000 ;
			15'h00001CA2 : data <= 8'b00000000 ;
			15'h00001CA3 : data <= 8'b00000000 ;
			15'h00001CA4 : data <= 8'b00000000 ;
			15'h00001CA5 : data <= 8'b00000000 ;
			15'h00001CA6 : data <= 8'b00000000 ;
			15'h00001CA7 : data <= 8'b00000000 ;
			15'h00001CA8 : data <= 8'b00000000 ;
			15'h00001CA9 : data <= 8'b00000000 ;
			15'h00001CAA : data <= 8'b00000000 ;
			15'h00001CAB : data <= 8'b00000000 ;
			15'h00001CAC : data <= 8'b00000000 ;
			15'h00001CAD : data <= 8'b00000000 ;
			15'h00001CAE : data <= 8'b00000000 ;
			15'h00001CAF : data <= 8'b00000000 ;
			15'h00001CB0 : data <= 8'b00000000 ;
			15'h00001CB1 : data <= 8'b00000000 ;
			15'h00001CB2 : data <= 8'b00000000 ;
			15'h00001CB3 : data <= 8'b00000000 ;
			15'h00001CB4 : data <= 8'b00000000 ;
			15'h00001CB5 : data <= 8'b00000000 ;
			15'h00001CB6 : data <= 8'b00000000 ;
			15'h00001CB7 : data <= 8'b00000000 ;
			15'h00001CB8 : data <= 8'b00000000 ;
			15'h00001CB9 : data <= 8'b00000000 ;
			15'h00001CBA : data <= 8'b00000000 ;
			15'h00001CBB : data <= 8'b00000000 ;
			15'h00001CBC : data <= 8'b00000000 ;
			15'h00001CBD : data <= 8'b00000000 ;
			15'h00001CBE : data <= 8'b00000000 ;
			15'h00001CBF : data <= 8'b00000000 ;
			15'h00001CC0 : data <= 8'b00000000 ;
			15'h00001CC1 : data <= 8'b00000000 ;
			15'h00001CC2 : data <= 8'b00000000 ;
			15'h00001CC3 : data <= 8'b00000000 ;
			15'h00001CC4 : data <= 8'b00000000 ;
			15'h00001CC5 : data <= 8'b00000000 ;
			15'h00001CC6 : data <= 8'b00000000 ;
			15'h00001CC7 : data <= 8'b00000000 ;
			15'h00001CC8 : data <= 8'b00000000 ;
			15'h00001CC9 : data <= 8'b00000000 ;
			15'h00001CCA : data <= 8'b00000000 ;
			15'h00001CCB : data <= 8'b00000000 ;
			15'h00001CCC : data <= 8'b00000000 ;
			15'h00001CCD : data <= 8'b00000000 ;
			15'h00001CCE : data <= 8'b00000000 ;
			15'h00001CCF : data <= 8'b00000000 ;
			15'h00001CD0 : data <= 8'b00000000 ;
			15'h00001CD1 : data <= 8'b00000000 ;
			15'h00001CD2 : data <= 8'b00000000 ;
			15'h00001CD3 : data <= 8'b00000000 ;
			15'h00001CD4 : data <= 8'b00000000 ;
			15'h00001CD5 : data <= 8'b00000000 ;
			15'h00001CD6 : data <= 8'b00000000 ;
			15'h00001CD7 : data <= 8'b00000000 ;
			15'h00001CD8 : data <= 8'b00000000 ;
			15'h00001CD9 : data <= 8'b00000000 ;
			15'h00001CDA : data <= 8'b00000000 ;
			15'h00001CDB : data <= 8'b00000000 ;
			15'h00001CDC : data <= 8'b00000000 ;
			15'h00001CDD : data <= 8'b00000000 ;
			15'h00001CDE : data <= 8'b00000000 ;
			15'h00001CDF : data <= 8'b00000000 ;
			15'h00001CE0 : data <= 8'b00000000 ;
			15'h00001CE1 : data <= 8'b00000000 ;
			15'h00001CE2 : data <= 8'b00000000 ;
			15'h00001CE3 : data <= 8'b00000000 ;
			15'h00001CE4 : data <= 8'b00000000 ;
			15'h00001CE5 : data <= 8'b00000000 ;
			15'h00001CE6 : data <= 8'b00000000 ;
			15'h00001CE7 : data <= 8'b00000000 ;
			15'h00001CE8 : data <= 8'b00000000 ;
			15'h00001CE9 : data <= 8'b00000000 ;
			15'h00001CEA : data <= 8'b00000000 ;
			15'h00001CEB : data <= 8'b00000000 ;
			15'h00001CEC : data <= 8'b00000000 ;
			15'h00001CED : data <= 8'b00000000 ;
			15'h00001CEE : data <= 8'b00000000 ;
			15'h00001CEF : data <= 8'b00000000 ;
			15'h00001CF0 : data <= 8'b00000000 ;
			15'h00001CF1 : data <= 8'b00000000 ;
			15'h00001CF2 : data <= 8'b00000000 ;
			15'h00001CF3 : data <= 8'b00000000 ;
			15'h00001CF4 : data <= 8'b00000000 ;
			15'h00001CF5 : data <= 8'b00000000 ;
			15'h00001CF6 : data <= 8'b00000000 ;
			15'h00001CF7 : data <= 8'b00000000 ;
			15'h00001CF8 : data <= 8'b00000000 ;
			15'h00001CF9 : data <= 8'b00000000 ;
			15'h00001CFA : data <= 8'b00000000 ;
			15'h00001CFB : data <= 8'b00000000 ;
			15'h00001CFC : data <= 8'b00000000 ;
			15'h00001CFD : data <= 8'b00000000 ;
			15'h00001CFE : data <= 8'b00000000 ;
			15'h00001CFF : data <= 8'b00000000 ;
			15'h00001D00 : data <= 8'b00000000 ;
			15'h00001D01 : data <= 8'b00000000 ;
			15'h00001D02 : data <= 8'b00000000 ;
			15'h00001D03 : data <= 8'b00000000 ;
			15'h00001D04 : data <= 8'b00000000 ;
			15'h00001D05 : data <= 8'b00000000 ;
			15'h00001D06 : data <= 8'b00000000 ;
			15'h00001D07 : data <= 8'b00000000 ;
			15'h00001D08 : data <= 8'b00000000 ;
			15'h00001D09 : data <= 8'b00000000 ;
			15'h00001D0A : data <= 8'b00000000 ;
			15'h00001D0B : data <= 8'b00000000 ;
			15'h00001D0C : data <= 8'b00000000 ;
			15'h00001D0D : data <= 8'b00000000 ;
			15'h00001D0E : data <= 8'b00000000 ;
			15'h00001D0F : data <= 8'b00000000 ;
			15'h00001D10 : data <= 8'b00000000 ;
			15'h00001D11 : data <= 8'b00000000 ;
			15'h00001D12 : data <= 8'b00000000 ;
			15'h00001D13 : data <= 8'b00000000 ;
			15'h00001D14 : data <= 8'b00000000 ;
			15'h00001D15 : data <= 8'b00000000 ;
			15'h00001D16 : data <= 8'b00000000 ;
			15'h00001D17 : data <= 8'b00000000 ;
			15'h00001D18 : data <= 8'b00000000 ;
			15'h00001D19 : data <= 8'b00000000 ;
			15'h00001D1A : data <= 8'b00000000 ;
			15'h00001D1B : data <= 8'b00000000 ;
			15'h00001D1C : data <= 8'b00000000 ;
			15'h00001D1D : data <= 8'b00000000 ;
			15'h00001D1E : data <= 8'b00000000 ;
			15'h00001D1F : data <= 8'b00000000 ;
			15'h00001D20 : data <= 8'b00000000 ;
			15'h00001D21 : data <= 8'b00000000 ;
			15'h00001D22 : data <= 8'b00000000 ;
			15'h00001D23 : data <= 8'b00000000 ;
			15'h00001D24 : data <= 8'b00000000 ;
			15'h00001D25 : data <= 8'b00000000 ;
			15'h00001D26 : data <= 8'b00000000 ;
			15'h00001D27 : data <= 8'b00000000 ;
			15'h00001D28 : data <= 8'b00000000 ;
			15'h00001D29 : data <= 8'b00000000 ;
			15'h00001D2A : data <= 8'b00000000 ;
			15'h00001D2B : data <= 8'b00000000 ;
			15'h00001D2C : data <= 8'b00000000 ;
			15'h00001D2D : data <= 8'b00000000 ;
			15'h00001D2E : data <= 8'b00000000 ;
			15'h00001D2F : data <= 8'b00000000 ;
			15'h00001D30 : data <= 8'b00000000 ;
			15'h00001D31 : data <= 8'b00000000 ;
			15'h00001D32 : data <= 8'b00000000 ;
			15'h00001D33 : data <= 8'b00000000 ;
			15'h00001D34 : data <= 8'b00000000 ;
			15'h00001D35 : data <= 8'b00000000 ;
			15'h00001D36 : data <= 8'b00000000 ;
			15'h00001D37 : data <= 8'b00000000 ;
			15'h00001D38 : data <= 8'b00000000 ;
			15'h00001D39 : data <= 8'b00000000 ;
			15'h00001D3A : data <= 8'b00000000 ;
			15'h00001D3B : data <= 8'b00000000 ;
			15'h00001D3C : data <= 8'b00000000 ;
			15'h00001D3D : data <= 8'b00000000 ;
			15'h00001D3E : data <= 8'b00000000 ;
			15'h00001D3F : data <= 8'b00000000 ;
			15'h00001D40 : data <= 8'b00000000 ;
			15'h00001D41 : data <= 8'b00000000 ;
			15'h00001D42 : data <= 8'b00000000 ;
			15'h00001D43 : data <= 8'b00000000 ;
			15'h00001D44 : data <= 8'b00000000 ;
			15'h00001D45 : data <= 8'b00000000 ;
			15'h00001D46 : data <= 8'b00000000 ;
			15'h00001D47 : data <= 8'b00000000 ;
			15'h00001D48 : data <= 8'b00000000 ;
			15'h00001D49 : data <= 8'b00000000 ;
			15'h00001D4A : data <= 8'b00000000 ;
			15'h00001D4B : data <= 8'b00000000 ;
			15'h00001D4C : data <= 8'b00000000 ;
			15'h00001D4D : data <= 8'b00000000 ;
			15'h00001D4E : data <= 8'b00000000 ;
			15'h00001D4F : data <= 8'b00000000 ;
			15'h00001D50 : data <= 8'b00000000 ;
			15'h00001D51 : data <= 8'b00000000 ;
			15'h00001D52 : data <= 8'b00000000 ;
			15'h00001D53 : data <= 8'b00000000 ;
			15'h00001D54 : data <= 8'b00000000 ;
			15'h00001D55 : data <= 8'b00000000 ;
			15'h00001D56 : data <= 8'b00000000 ;
			15'h00001D57 : data <= 8'b00000000 ;
			15'h00001D58 : data <= 8'b00000000 ;
			15'h00001D59 : data <= 8'b00000000 ;
			15'h00001D5A : data <= 8'b00000000 ;
			15'h00001D5B : data <= 8'b00000000 ;
			15'h00001D5C : data <= 8'b00000000 ;
			15'h00001D5D : data <= 8'b00000000 ;
			15'h00001D5E : data <= 8'b00000000 ;
			15'h00001D5F : data <= 8'b00000000 ;
			15'h00001D60 : data <= 8'b00000000 ;
			15'h00001D61 : data <= 8'b00000000 ;
			15'h00001D62 : data <= 8'b00000000 ;
			15'h00001D63 : data <= 8'b00000000 ;
			15'h00001D64 : data <= 8'b00000000 ;
			15'h00001D65 : data <= 8'b00000000 ;
			15'h00001D66 : data <= 8'b00000000 ;
			15'h00001D67 : data <= 8'b00000000 ;
			15'h00001D68 : data <= 8'b00000000 ;
			15'h00001D69 : data <= 8'b00000000 ;
			15'h00001D6A : data <= 8'b00000000 ;
			15'h00001D6B : data <= 8'b00000000 ;
			15'h00001D6C : data <= 8'b00000000 ;
			15'h00001D6D : data <= 8'b00000000 ;
			15'h00001D6E : data <= 8'b00000000 ;
			15'h00001D6F : data <= 8'b00000000 ;
			15'h00001D70 : data <= 8'b00000000 ;
			15'h00001D71 : data <= 8'b00000000 ;
			15'h00001D72 : data <= 8'b00000000 ;
			15'h00001D73 : data <= 8'b00000000 ;
			15'h00001D74 : data <= 8'b00000000 ;
			15'h00001D75 : data <= 8'b00000000 ;
			15'h00001D76 : data <= 8'b00000000 ;
			15'h00001D77 : data <= 8'b00000000 ;
			15'h00001D78 : data <= 8'b00000000 ;
			15'h00001D79 : data <= 8'b00000000 ;
			15'h00001D7A : data <= 8'b00000000 ;
			15'h00001D7B : data <= 8'b00000000 ;
			15'h00001D7C : data <= 8'b00000000 ;
			15'h00001D7D : data <= 8'b00000000 ;
			15'h00001D7E : data <= 8'b00000000 ;
			15'h00001D7F : data <= 8'b00000000 ;
			15'h00001D80 : data <= 8'b00000000 ;
			15'h00001D81 : data <= 8'b00000000 ;
			15'h00001D82 : data <= 8'b00000000 ;
			15'h00001D83 : data <= 8'b00000000 ;
			15'h00001D84 : data <= 8'b00000000 ;
			15'h00001D85 : data <= 8'b00000000 ;
			15'h00001D86 : data <= 8'b00000000 ;
			15'h00001D87 : data <= 8'b00000000 ;
			15'h00001D88 : data <= 8'b00000000 ;
			15'h00001D89 : data <= 8'b00000000 ;
			15'h00001D8A : data <= 8'b00000000 ;
			15'h00001D8B : data <= 8'b00000000 ;
			15'h00001D8C : data <= 8'b00000000 ;
			15'h00001D8D : data <= 8'b00000000 ;
			15'h00001D8E : data <= 8'b00000000 ;
			15'h00001D8F : data <= 8'b00000000 ;
			15'h00001D90 : data <= 8'b00000000 ;
			15'h00001D91 : data <= 8'b00000000 ;
			15'h00001D92 : data <= 8'b00000000 ;
			15'h00001D93 : data <= 8'b00000000 ;
			15'h00001D94 : data <= 8'b00000000 ;
			15'h00001D95 : data <= 8'b00000000 ;
			15'h00001D96 : data <= 8'b00000000 ;
			15'h00001D97 : data <= 8'b00000000 ;
			15'h00001D98 : data <= 8'b00000000 ;
			15'h00001D99 : data <= 8'b00000000 ;
			15'h00001D9A : data <= 8'b00000000 ;
			15'h00001D9B : data <= 8'b00000000 ;
			15'h00001D9C : data <= 8'b00000000 ;
			15'h00001D9D : data <= 8'b00000000 ;
			15'h00001D9E : data <= 8'b00000000 ;
			15'h00001D9F : data <= 8'b00000000 ;
			15'h00001DA0 : data <= 8'b00000000 ;
			15'h00001DA1 : data <= 8'b00000000 ;
			15'h00001DA2 : data <= 8'b00000000 ;
			15'h00001DA3 : data <= 8'b00000000 ;
			15'h00001DA4 : data <= 8'b00000000 ;
			15'h00001DA5 : data <= 8'b00000000 ;
			15'h00001DA6 : data <= 8'b00000000 ;
			15'h00001DA7 : data <= 8'b00000000 ;
			15'h00001DA8 : data <= 8'b00000000 ;
			15'h00001DA9 : data <= 8'b00000000 ;
			15'h00001DAA : data <= 8'b00000000 ;
			15'h00001DAB : data <= 8'b00000000 ;
			15'h00001DAC : data <= 8'b00000000 ;
			15'h00001DAD : data <= 8'b00000000 ;
			15'h00001DAE : data <= 8'b00000000 ;
			15'h00001DAF : data <= 8'b00000000 ;
			15'h00001DB0 : data <= 8'b00000000 ;
			15'h00001DB1 : data <= 8'b00000000 ;
			15'h00001DB2 : data <= 8'b00000000 ;
			15'h00001DB3 : data <= 8'b00000000 ;
			15'h00001DB4 : data <= 8'b00000000 ;
			15'h00001DB5 : data <= 8'b00000000 ;
			15'h00001DB6 : data <= 8'b00000000 ;
			15'h00001DB7 : data <= 8'b00000000 ;
			15'h00001DB8 : data <= 8'b00000000 ;
			15'h00001DB9 : data <= 8'b00000000 ;
			15'h00001DBA : data <= 8'b00000000 ;
			15'h00001DBB : data <= 8'b00000000 ;
			15'h00001DBC : data <= 8'b00000000 ;
			15'h00001DBD : data <= 8'b00000000 ;
			15'h00001DBE : data <= 8'b00000000 ;
			15'h00001DBF : data <= 8'b00000000 ;
			15'h00001DC0 : data <= 8'b00000000 ;
			15'h00001DC1 : data <= 8'b00000000 ;
			15'h00001DC2 : data <= 8'b00000000 ;
			15'h00001DC3 : data <= 8'b00000000 ;
			15'h00001DC4 : data <= 8'b00000000 ;
			15'h00001DC5 : data <= 8'b00000000 ;
			15'h00001DC6 : data <= 8'b00000000 ;
			15'h00001DC7 : data <= 8'b00000000 ;
			15'h00001DC8 : data <= 8'b00000000 ;
			15'h00001DC9 : data <= 8'b00000000 ;
			15'h00001DCA : data <= 8'b00000000 ;
			15'h00001DCB : data <= 8'b00000000 ;
			15'h00001DCC : data <= 8'b00000000 ;
			15'h00001DCD : data <= 8'b00000000 ;
			15'h00001DCE : data <= 8'b00000000 ;
			15'h00001DCF : data <= 8'b00000000 ;
			15'h00001DD0 : data <= 8'b00000000 ;
			15'h00001DD1 : data <= 8'b00000000 ;
			15'h00001DD2 : data <= 8'b00000000 ;
			15'h00001DD3 : data <= 8'b00000000 ;
			15'h00001DD4 : data <= 8'b00000000 ;
			15'h00001DD5 : data <= 8'b00000000 ;
			15'h00001DD6 : data <= 8'b00000000 ;
			15'h00001DD7 : data <= 8'b00000000 ;
			15'h00001DD8 : data <= 8'b00000000 ;
			15'h00001DD9 : data <= 8'b00000000 ;
			15'h00001DDA : data <= 8'b00000000 ;
			15'h00001DDB : data <= 8'b00000000 ;
			15'h00001DDC : data <= 8'b00000000 ;
			15'h00001DDD : data <= 8'b00000000 ;
			15'h00001DDE : data <= 8'b00000000 ;
			15'h00001DDF : data <= 8'b00000000 ;
			15'h00001DE0 : data <= 8'b00000000 ;
			15'h00001DE1 : data <= 8'b00000000 ;
			15'h00001DE2 : data <= 8'b00000000 ;
			15'h00001DE3 : data <= 8'b00000000 ;
			15'h00001DE4 : data <= 8'b00000000 ;
			15'h00001DE5 : data <= 8'b00000000 ;
			15'h00001DE6 : data <= 8'b00000000 ;
			15'h00001DE7 : data <= 8'b00000000 ;
			15'h00001DE8 : data <= 8'b00000000 ;
			15'h00001DE9 : data <= 8'b00000000 ;
			15'h00001DEA : data <= 8'b00000000 ;
			15'h00001DEB : data <= 8'b00000000 ;
			15'h00001DEC : data <= 8'b00000000 ;
			15'h00001DED : data <= 8'b00000000 ;
			15'h00001DEE : data <= 8'b00000000 ;
			15'h00001DEF : data <= 8'b00000000 ;
			15'h00001DF0 : data <= 8'b00000000 ;
			15'h00001DF1 : data <= 8'b00000000 ;
			15'h00001DF2 : data <= 8'b00000000 ;
			15'h00001DF3 : data <= 8'b00000000 ;
			15'h00001DF4 : data <= 8'b00000000 ;
			15'h00001DF5 : data <= 8'b00000000 ;
			15'h00001DF6 : data <= 8'b00000000 ;
			15'h00001DF7 : data <= 8'b00000000 ;
			15'h00001DF8 : data <= 8'b00000000 ;
			15'h00001DF9 : data <= 8'b00000000 ;
			15'h00001DFA : data <= 8'b00000000 ;
			15'h00001DFB : data <= 8'b00000000 ;
			15'h00001DFC : data <= 8'b00000000 ;
			15'h00001DFD : data <= 8'b00000000 ;
			15'h00001DFE : data <= 8'b00000000 ;
			15'h00001DFF : data <= 8'b00000000 ;
			15'h00001E00 : data <= 8'b00000000 ;
			15'h00001E01 : data <= 8'b00000000 ;
			15'h00001E02 : data <= 8'b00000000 ;
			15'h00001E03 : data <= 8'b00000000 ;
			15'h00001E04 : data <= 8'b00000000 ;
			15'h00001E05 : data <= 8'b00000000 ;
			15'h00001E06 : data <= 8'b00000000 ;
			15'h00001E07 : data <= 8'b00000000 ;
			15'h00001E08 : data <= 8'b00000000 ;
			15'h00001E09 : data <= 8'b00000000 ;
			15'h00001E0A : data <= 8'b00000000 ;
			15'h00001E0B : data <= 8'b00000000 ;
			15'h00001E0C : data <= 8'b00000000 ;
			15'h00001E0D : data <= 8'b00000000 ;
			15'h00001E0E : data <= 8'b00000000 ;
			15'h00001E0F : data <= 8'b00000000 ;
			15'h00001E10 : data <= 8'b00000000 ;
			15'h00001E11 : data <= 8'b00000000 ;
			15'h00001E12 : data <= 8'b00000000 ;
			15'h00001E13 : data <= 8'b00000000 ;
			15'h00001E14 : data <= 8'b00000000 ;
			15'h00001E15 : data <= 8'b00000000 ;
			15'h00001E16 : data <= 8'b00000000 ;
			15'h00001E17 : data <= 8'b00000000 ;
			15'h00001E18 : data <= 8'b00000000 ;
			15'h00001E19 : data <= 8'b00000000 ;
			15'h00001E1A : data <= 8'b00000000 ;
			15'h00001E1B : data <= 8'b00000000 ;
			15'h00001E1C : data <= 8'b00000000 ;
			15'h00001E1D : data <= 8'b00000000 ;
			15'h00001E1E : data <= 8'b00000000 ;
			15'h00001E1F : data <= 8'b00000000 ;
			15'h00001E20 : data <= 8'b00000000 ;
			15'h00001E21 : data <= 8'b00000000 ;
			15'h00001E22 : data <= 8'b00000000 ;
			15'h00001E23 : data <= 8'b00000000 ;
			15'h00001E24 : data <= 8'b00000000 ;
			15'h00001E25 : data <= 8'b00000000 ;
			15'h00001E26 : data <= 8'b00000000 ;
			15'h00001E27 : data <= 8'b00000000 ;
			15'h00001E28 : data <= 8'b00000000 ;
			15'h00001E29 : data <= 8'b00000000 ;
			15'h00001E2A : data <= 8'b00000000 ;
			15'h00001E2B : data <= 8'b00000000 ;
			15'h00001E2C : data <= 8'b00000000 ;
			15'h00001E2D : data <= 8'b00000000 ;
			15'h00001E2E : data <= 8'b00000000 ;
			15'h00001E2F : data <= 8'b00000000 ;
			15'h00001E30 : data <= 8'b00000000 ;
			15'h00001E31 : data <= 8'b00000000 ;
			15'h00001E32 : data <= 8'b00000000 ;
			15'h00001E33 : data <= 8'b00000000 ;
			15'h00001E34 : data <= 8'b00000000 ;
			15'h00001E35 : data <= 8'b00000000 ;
			15'h00001E36 : data <= 8'b00000000 ;
			15'h00001E37 : data <= 8'b00000000 ;
			15'h00001E38 : data <= 8'b00000000 ;
			15'h00001E39 : data <= 8'b00000000 ;
			15'h00001E3A : data <= 8'b00000000 ;
			15'h00001E3B : data <= 8'b00000000 ;
			15'h00001E3C : data <= 8'b00000000 ;
			15'h00001E3D : data <= 8'b00000000 ;
			15'h00001E3E : data <= 8'b00000000 ;
			15'h00001E3F : data <= 8'b00000000 ;
			15'h00001E40 : data <= 8'b00000000 ;
			15'h00001E41 : data <= 8'b00000000 ;
			15'h00001E42 : data <= 8'b00000000 ;
			15'h00001E43 : data <= 8'b00000000 ;
			15'h00001E44 : data <= 8'b00000000 ;
			15'h00001E45 : data <= 8'b00000000 ;
			15'h00001E46 : data <= 8'b00000000 ;
			15'h00001E47 : data <= 8'b00000000 ;
			15'h00001E48 : data <= 8'b00000000 ;
			15'h00001E49 : data <= 8'b00000000 ;
			15'h00001E4A : data <= 8'b00000000 ;
			15'h00001E4B : data <= 8'b00000000 ;
			15'h00001E4C : data <= 8'b00000000 ;
			15'h00001E4D : data <= 8'b00000000 ;
			15'h00001E4E : data <= 8'b00000000 ;
			15'h00001E4F : data <= 8'b00000000 ;
			15'h00001E50 : data <= 8'b00000000 ;
			15'h00001E51 : data <= 8'b00000000 ;
			15'h00001E52 : data <= 8'b00000000 ;
			15'h00001E53 : data <= 8'b00000000 ;
			15'h00001E54 : data <= 8'b00000000 ;
			15'h00001E55 : data <= 8'b00000000 ;
			15'h00001E56 : data <= 8'b00000000 ;
			15'h00001E57 : data <= 8'b00000000 ;
			15'h00001E58 : data <= 8'b00000000 ;
			15'h00001E59 : data <= 8'b00000000 ;
			15'h00001E5A : data <= 8'b00000000 ;
			15'h00001E5B : data <= 8'b00000000 ;
			15'h00001E5C : data <= 8'b00000000 ;
			15'h00001E5D : data <= 8'b00000000 ;
			15'h00001E5E : data <= 8'b00000000 ;
			15'h00001E5F : data <= 8'b00000000 ;
			15'h00001E60 : data <= 8'b00000000 ;
			15'h00001E61 : data <= 8'b00000000 ;
			15'h00001E62 : data <= 8'b00000000 ;
			15'h00001E63 : data <= 8'b00000000 ;
			15'h00001E64 : data <= 8'b00000000 ;
			15'h00001E65 : data <= 8'b00000000 ;
			15'h00001E66 : data <= 8'b00000000 ;
			15'h00001E67 : data <= 8'b00000000 ;
			15'h00001E68 : data <= 8'b00000000 ;
			15'h00001E69 : data <= 8'b00000000 ;
			15'h00001E6A : data <= 8'b00000000 ;
			15'h00001E6B : data <= 8'b00000000 ;
			15'h00001E6C : data <= 8'b00000000 ;
			15'h00001E6D : data <= 8'b00000000 ;
			15'h00001E6E : data <= 8'b00000000 ;
			15'h00001E6F : data <= 8'b00000000 ;
			15'h00001E70 : data <= 8'b00000000 ;
			15'h00001E71 : data <= 8'b00000000 ;
			15'h00001E72 : data <= 8'b00000000 ;
			15'h00001E73 : data <= 8'b00000000 ;
			15'h00001E74 : data <= 8'b00000000 ;
			15'h00001E75 : data <= 8'b00000000 ;
			15'h00001E76 : data <= 8'b00000000 ;
			15'h00001E77 : data <= 8'b00000000 ;
			15'h00001E78 : data <= 8'b00000000 ;
			15'h00001E79 : data <= 8'b00000000 ;
			15'h00001E7A : data <= 8'b00000000 ;
			15'h00001E7B : data <= 8'b00000000 ;
			15'h00001E7C : data <= 8'b00000000 ;
			15'h00001E7D : data <= 8'b00000000 ;
			15'h00001E7E : data <= 8'b00000000 ;
			15'h00001E7F : data <= 8'b00000000 ;
			15'h00001E80 : data <= 8'b00000000 ;
			15'h00001E81 : data <= 8'b00000000 ;
			15'h00001E82 : data <= 8'b00000000 ;
			15'h00001E83 : data <= 8'b00000000 ;
			15'h00001E84 : data <= 8'b00000000 ;
			15'h00001E85 : data <= 8'b00000000 ;
			15'h00001E86 : data <= 8'b00000000 ;
			15'h00001E87 : data <= 8'b00000000 ;
			15'h00001E88 : data <= 8'b00000000 ;
			15'h00001E89 : data <= 8'b00000000 ;
			15'h00001E8A : data <= 8'b00000000 ;
			15'h00001E8B : data <= 8'b00000000 ;
			15'h00001E8C : data <= 8'b00000000 ;
			15'h00001E8D : data <= 8'b00000000 ;
			15'h00001E8E : data <= 8'b00000000 ;
			15'h00001E8F : data <= 8'b00000000 ;
			15'h00001E90 : data <= 8'b00000000 ;
			15'h00001E91 : data <= 8'b00000000 ;
			15'h00001E92 : data <= 8'b00000000 ;
			15'h00001E93 : data <= 8'b00000000 ;
			15'h00001E94 : data <= 8'b00000000 ;
			15'h00001E95 : data <= 8'b00000000 ;
			15'h00001E96 : data <= 8'b00000000 ;
			15'h00001E97 : data <= 8'b00000000 ;
			15'h00001E98 : data <= 8'b00000000 ;
			15'h00001E99 : data <= 8'b00000000 ;
			15'h00001E9A : data <= 8'b00000000 ;
			15'h00001E9B : data <= 8'b00000000 ;
			15'h00001E9C : data <= 8'b00000000 ;
			15'h00001E9D : data <= 8'b00000000 ;
			15'h00001E9E : data <= 8'b00000000 ;
			15'h00001E9F : data <= 8'b00000000 ;
			15'h00001EA0 : data <= 8'b00000000 ;
			15'h00001EA1 : data <= 8'b00000000 ;
			15'h00001EA2 : data <= 8'b00000000 ;
			15'h00001EA3 : data <= 8'b00000000 ;
			15'h00001EA4 : data <= 8'b00000000 ;
			15'h00001EA5 : data <= 8'b00000000 ;
			15'h00001EA6 : data <= 8'b00000000 ;
			15'h00001EA7 : data <= 8'b00000000 ;
			15'h00001EA8 : data <= 8'b00000000 ;
			15'h00001EA9 : data <= 8'b00000000 ;
			15'h00001EAA : data <= 8'b00000000 ;
			15'h00001EAB : data <= 8'b00000000 ;
			15'h00001EAC : data <= 8'b00000000 ;
			15'h00001EAD : data <= 8'b00000000 ;
			15'h00001EAE : data <= 8'b00000000 ;
			15'h00001EAF : data <= 8'b00000000 ;
			15'h00001EB0 : data <= 8'b00000000 ;
			15'h00001EB1 : data <= 8'b00000000 ;
			15'h00001EB2 : data <= 8'b00000000 ;
			15'h00001EB3 : data <= 8'b00000000 ;
			15'h00001EB4 : data <= 8'b00000000 ;
			15'h00001EB5 : data <= 8'b00000000 ;
			15'h00001EB6 : data <= 8'b00000000 ;
			15'h00001EB7 : data <= 8'b00000000 ;
			15'h00001EB8 : data <= 8'b00000000 ;
			15'h00001EB9 : data <= 8'b00000000 ;
			15'h00001EBA : data <= 8'b00000000 ;
			15'h00001EBB : data <= 8'b00000000 ;
			15'h00001EBC : data <= 8'b00000000 ;
			15'h00001EBD : data <= 8'b00000000 ;
			15'h00001EBE : data <= 8'b00000000 ;
			15'h00001EBF : data <= 8'b00000000 ;
			15'h00001EC0 : data <= 8'b00000000 ;
			15'h00001EC1 : data <= 8'b00000000 ;
			15'h00001EC2 : data <= 8'b00000000 ;
			15'h00001EC3 : data <= 8'b00000000 ;
			15'h00001EC4 : data <= 8'b00000000 ;
			15'h00001EC5 : data <= 8'b00000000 ;
			15'h00001EC6 : data <= 8'b00000000 ;
			15'h00001EC7 : data <= 8'b00000000 ;
			15'h00001EC8 : data <= 8'b00000000 ;
			15'h00001EC9 : data <= 8'b00000000 ;
			15'h00001ECA : data <= 8'b00000000 ;
			15'h00001ECB : data <= 8'b00000000 ;
			15'h00001ECC : data <= 8'b00000000 ;
			15'h00001ECD : data <= 8'b00000000 ;
			15'h00001ECE : data <= 8'b00000000 ;
			15'h00001ECF : data <= 8'b00000000 ;
			15'h00001ED0 : data <= 8'b00000000 ;
			15'h00001ED1 : data <= 8'b00000000 ;
			15'h00001ED2 : data <= 8'b00000000 ;
			15'h00001ED3 : data <= 8'b00000000 ;
			15'h00001ED4 : data <= 8'b00000000 ;
			15'h00001ED5 : data <= 8'b00000000 ;
			15'h00001ED6 : data <= 8'b00000000 ;
			15'h00001ED7 : data <= 8'b00000000 ;
			15'h00001ED8 : data <= 8'b00000000 ;
			15'h00001ED9 : data <= 8'b00000000 ;
			15'h00001EDA : data <= 8'b00000000 ;
			15'h00001EDB : data <= 8'b00000000 ;
			15'h00001EDC : data <= 8'b00000000 ;
			15'h00001EDD : data <= 8'b00000000 ;
			15'h00001EDE : data <= 8'b00000000 ;
			15'h00001EDF : data <= 8'b00000000 ;
			15'h00001EE0 : data <= 8'b00000000 ;
			15'h00001EE1 : data <= 8'b00000000 ;
			15'h00001EE2 : data <= 8'b00000000 ;
			15'h00001EE3 : data <= 8'b00000000 ;
			15'h00001EE4 : data <= 8'b00000000 ;
			15'h00001EE5 : data <= 8'b00000000 ;
			15'h00001EE6 : data <= 8'b00000000 ;
			15'h00001EE7 : data <= 8'b00000000 ;
			15'h00001EE8 : data <= 8'b00000000 ;
			15'h00001EE9 : data <= 8'b00000000 ;
			15'h00001EEA : data <= 8'b00000000 ;
			15'h00001EEB : data <= 8'b00000000 ;
			15'h00001EEC : data <= 8'b00000000 ;
			15'h00001EED : data <= 8'b00000000 ;
			15'h00001EEE : data <= 8'b00000000 ;
			15'h00001EEF : data <= 8'b00000000 ;
			15'h00001EF0 : data <= 8'b00000000 ;
			15'h00001EF1 : data <= 8'b00000000 ;
			15'h00001EF2 : data <= 8'b00000000 ;
			15'h00001EF3 : data <= 8'b00000000 ;
			15'h00001EF4 : data <= 8'b00000000 ;
			15'h00001EF5 : data <= 8'b00000000 ;
			15'h00001EF6 : data <= 8'b00000000 ;
			15'h00001EF7 : data <= 8'b00000000 ;
			15'h00001EF8 : data <= 8'b00000000 ;
			15'h00001EF9 : data <= 8'b00000000 ;
			15'h00001EFA : data <= 8'b00000000 ;
			15'h00001EFB : data <= 8'b00000000 ;
			15'h00001EFC : data <= 8'b00000000 ;
			15'h00001EFD : data <= 8'b00000000 ;
			15'h00001EFE : data <= 8'b00000000 ;
			15'h00001EFF : data <= 8'b00000000 ;
			15'h00001F00 : data <= 8'b00000000 ;
			15'h00001F01 : data <= 8'b00000000 ;
			15'h00001F02 : data <= 8'b00000000 ;
			15'h00001F03 : data <= 8'b00000000 ;
			15'h00001F04 : data <= 8'b00000000 ;
			15'h00001F05 : data <= 8'b00000000 ;
			15'h00001F06 : data <= 8'b00000000 ;
			15'h00001F07 : data <= 8'b00000000 ;
			15'h00001F08 : data <= 8'b00000000 ;
			15'h00001F09 : data <= 8'b00000000 ;
			15'h00001F0A : data <= 8'b00000000 ;
			15'h00001F0B : data <= 8'b00000000 ;
			15'h00001F0C : data <= 8'b00000000 ;
			15'h00001F0D : data <= 8'b00000000 ;
			15'h00001F0E : data <= 8'b00000000 ;
			15'h00001F0F : data <= 8'b00000000 ;
			15'h00001F10 : data <= 8'b00000000 ;
			15'h00001F11 : data <= 8'b00000000 ;
			15'h00001F12 : data <= 8'b00000000 ;
			15'h00001F13 : data <= 8'b00000000 ;
			15'h00001F14 : data <= 8'b00000000 ;
			15'h00001F15 : data <= 8'b00000000 ;
			15'h00001F16 : data <= 8'b00000000 ;
			15'h00001F17 : data <= 8'b00000000 ;
			15'h00001F18 : data <= 8'b00000000 ;
			15'h00001F19 : data <= 8'b00000000 ;
			15'h00001F1A : data <= 8'b00000000 ;
			15'h00001F1B : data <= 8'b00000000 ;
			15'h00001F1C : data <= 8'b00000000 ;
			15'h00001F1D : data <= 8'b00000000 ;
			15'h00001F1E : data <= 8'b00000000 ;
			15'h00001F1F : data <= 8'b00000000 ;
			15'h00001F20 : data <= 8'b00000000 ;
			15'h00001F21 : data <= 8'b00000000 ;
			15'h00001F22 : data <= 8'b00000000 ;
			15'h00001F23 : data <= 8'b00000000 ;
			15'h00001F24 : data <= 8'b00000000 ;
			15'h00001F25 : data <= 8'b00000000 ;
			15'h00001F26 : data <= 8'b00000000 ;
			15'h00001F27 : data <= 8'b00000000 ;
			15'h00001F28 : data <= 8'b00000000 ;
			15'h00001F29 : data <= 8'b00000000 ;
			15'h00001F2A : data <= 8'b00000000 ;
			15'h00001F2B : data <= 8'b00000000 ;
			15'h00001F2C : data <= 8'b00000000 ;
			15'h00001F2D : data <= 8'b00000000 ;
			15'h00001F2E : data <= 8'b00000000 ;
			15'h00001F2F : data <= 8'b00000000 ;
			15'h00001F30 : data <= 8'b00000000 ;
			15'h00001F31 : data <= 8'b00000000 ;
			15'h00001F32 : data <= 8'b00000000 ;
			15'h00001F33 : data <= 8'b00000000 ;
			15'h00001F34 : data <= 8'b00000000 ;
			15'h00001F35 : data <= 8'b00000000 ;
			15'h00001F36 : data <= 8'b00000000 ;
			15'h00001F37 : data <= 8'b00000000 ;
			15'h00001F38 : data <= 8'b00000000 ;
			15'h00001F39 : data <= 8'b00000000 ;
			15'h00001F3A : data <= 8'b00000000 ;
			15'h00001F3B : data <= 8'b00000000 ;
			15'h00001F3C : data <= 8'b00000000 ;
			15'h00001F3D : data <= 8'b00000000 ;
			15'h00001F3E : data <= 8'b00000000 ;
			15'h00001F3F : data <= 8'b00000000 ;
			15'h00001F40 : data <= 8'b00000000 ;
			15'h00001F41 : data <= 8'b00000000 ;
			15'h00001F42 : data <= 8'b00000000 ;
			15'h00001F43 : data <= 8'b00000000 ;
			15'h00001F44 : data <= 8'b00000000 ;
			15'h00001F45 : data <= 8'b00000000 ;
			15'h00001F46 : data <= 8'b00000000 ;
			15'h00001F47 : data <= 8'b00000000 ;
			15'h00001F48 : data <= 8'b00000000 ;
			15'h00001F49 : data <= 8'b00000000 ;
			15'h00001F4A : data <= 8'b00000000 ;
			15'h00001F4B : data <= 8'b00000000 ;
			15'h00001F4C : data <= 8'b00000000 ;
			15'h00001F4D : data <= 8'b00000000 ;
			15'h00001F4E : data <= 8'b00000000 ;
			15'h00001F4F : data <= 8'b00000000 ;
			15'h00001F50 : data <= 8'b00000000 ;
			15'h00001F51 : data <= 8'b00000000 ;
			15'h00001F52 : data <= 8'b00000000 ;
			15'h00001F53 : data <= 8'b00000000 ;
			15'h00001F54 : data <= 8'b00000000 ;
			15'h00001F55 : data <= 8'b00000000 ;
			15'h00001F56 : data <= 8'b00000000 ;
			15'h00001F57 : data <= 8'b00000000 ;
			15'h00001F58 : data <= 8'b00000000 ;
			15'h00001F59 : data <= 8'b00000000 ;
			15'h00001F5A : data <= 8'b00000000 ;
			15'h00001F5B : data <= 8'b00000000 ;
			15'h00001F5C : data <= 8'b00000000 ;
			15'h00001F5D : data <= 8'b00000000 ;
			15'h00001F5E : data <= 8'b00000000 ;
			15'h00001F5F : data <= 8'b00000000 ;
			15'h00001F60 : data <= 8'b00000000 ;
			15'h00001F61 : data <= 8'b00000000 ;
			15'h00001F62 : data <= 8'b00000000 ;
			15'h00001F63 : data <= 8'b00000000 ;
			15'h00001F64 : data <= 8'b00000000 ;
			15'h00001F65 : data <= 8'b00000000 ;
			15'h00001F66 : data <= 8'b00000000 ;
			15'h00001F67 : data <= 8'b00000000 ;
			15'h00001F68 : data <= 8'b00000000 ;
			15'h00001F69 : data <= 8'b00000000 ;
			15'h00001F6A : data <= 8'b00000000 ;
			15'h00001F6B : data <= 8'b00000000 ;
			15'h00001F6C : data <= 8'b00000000 ;
			15'h00001F6D : data <= 8'b00000000 ;
			15'h00001F6E : data <= 8'b00000000 ;
			15'h00001F6F : data <= 8'b00000000 ;
			15'h00001F70 : data <= 8'b00000000 ;
			15'h00001F71 : data <= 8'b00000000 ;
			15'h00001F72 : data <= 8'b00000000 ;
			15'h00001F73 : data <= 8'b00000000 ;
			15'h00001F74 : data <= 8'b00000000 ;
			15'h00001F75 : data <= 8'b00000000 ;
			15'h00001F76 : data <= 8'b00000000 ;
			15'h00001F77 : data <= 8'b00000000 ;
			15'h00001F78 : data <= 8'b00000000 ;
			15'h00001F79 : data <= 8'b00000000 ;
			15'h00001F7A : data <= 8'b00000000 ;
			15'h00001F7B : data <= 8'b00000000 ;
			15'h00001F7C : data <= 8'b00000000 ;
			15'h00001F7D : data <= 8'b00000000 ;
			15'h00001F7E : data <= 8'b00000000 ;
			15'h00001F7F : data <= 8'b00000000 ;
			15'h00001F80 : data <= 8'b00000000 ;
			15'h00001F81 : data <= 8'b00000000 ;
			15'h00001F82 : data <= 8'b00000000 ;
			15'h00001F83 : data <= 8'b00000000 ;
			15'h00001F84 : data <= 8'b00000000 ;
			15'h00001F85 : data <= 8'b00000000 ;
			15'h00001F86 : data <= 8'b00000000 ;
			15'h00001F87 : data <= 8'b00000000 ;
			15'h00001F88 : data <= 8'b00000000 ;
			15'h00001F89 : data <= 8'b00000000 ;
			15'h00001F8A : data <= 8'b00000000 ;
			15'h00001F8B : data <= 8'b00000000 ;
			15'h00001F8C : data <= 8'b00000000 ;
			15'h00001F8D : data <= 8'b00000000 ;
			15'h00001F8E : data <= 8'b00000000 ;
			15'h00001F8F : data <= 8'b00000000 ;
			15'h00001F90 : data <= 8'b00000000 ;
			15'h00001F91 : data <= 8'b00000000 ;
			15'h00001F92 : data <= 8'b00000000 ;
			15'h00001F93 : data <= 8'b00000000 ;
			15'h00001F94 : data <= 8'b00000000 ;
			15'h00001F95 : data <= 8'b00000000 ;
			15'h00001F96 : data <= 8'b00000000 ;
			15'h00001F97 : data <= 8'b00000000 ;
			15'h00001F98 : data <= 8'b00000000 ;
			15'h00001F99 : data <= 8'b00000000 ;
			15'h00001F9A : data <= 8'b00000000 ;
			15'h00001F9B : data <= 8'b00000000 ;
			15'h00001F9C : data <= 8'b00000000 ;
			15'h00001F9D : data <= 8'b00000000 ;
			15'h00001F9E : data <= 8'b00000000 ;
			15'h00001F9F : data <= 8'b00000000 ;
			15'h00001FA0 : data <= 8'b00000000 ;
			15'h00001FA1 : data <= 8'b00000000 ;
			15'h00001FA2 : data <= 8'b00000000 ;
			15'h00001FA3 : data <= 8'b00000000 ;
			15'h00001FA4 : data <= 8'b00000000 ;
			15'h00001FA5 : data <= 8'b00000000 ;
			15'h00001FA6 : data <= 8'b00000000 ;
			15'h00001FA7 : data <= 8'b00000000 ;
			15'h00001FA8 : data <= 8'b00000000 ;
			15'h00001FA9 : data <= 8'b00000000 ;
			15'h00001FAA : data <= 8'b00000000 ;
			15'h00001FAB : data <= 8'b00000000 ;
			15'h00001FAC : data <= 8'b00000000 ;
			15'h00001FAD : data <= 8'b00000000 ;
			15'h00001FAE : data <= 8'b00000000 ;
			15'h00001FAF : data <= 8'b00000000 ;
			15'h00001FB0 : data <= 8'b00000000 ;
			15'h00001FB1 : data <= 8'b00000000 ;
			15'h00001FB2 : data <= 8'b00000000 ;
			15'h00001FB3 : data <= 8'b00000000 ;
			15'h00001FB4 : data <= 8'b00000000 ;
			15'h00001FB5 : data <= 8'b00000000 ;
			15'h00001FB6 : data <= 8'b00000000 ;
			15'h00001FB7 : data <= 8'b00000000 ;
			15'h00001FB8 : data <= 8'b00000000 ;
			15'h00001FB9 : data <= 8'b00000000 ;
			15'h00001FBA : data <= 8'b00000000 ;
			15'h00001FBB : data <= 8'b00000000 ;
			15'h00001FBC : data <= 8'b00000000 ;
			15'h00001FBD : data <= 8'b00000000 ;
			15'h00001FBE : data <= 8'b00000000 ;
			15'h00001FBF : data <= 8'b00000000 ;
			15'h00001FC0 : data <= 8'b00000000 ;
			15'h00001FC1 : data <= 8'b00000000 ;
			15'h00001FC2 : data <= 8'b00000000 ;
			15'h00001FC3 : data <= 8'b00000000 ;
			15'h00001FC4 : data <= 8'b00000000 ;
			15'h00001FC5 : data <= 8'b00000000 ;
			15'h00001FC6 : data <= 8'b00000000 ;
			15'h00001FC7 : data <= 8'b00000000 ;
			15'h00001FC8 : data <= 8'b00000000 ;
			15'h00001FC9 : data <= 8'b00000000 ;
			15'h00001FCA : data <= 8'b00000000 ;
			15'h00001FCB : data <= 8'b00000000 ;
			15'h00001FCC : data <= 8'b00000000 ;
			15'h00001FCD : data <= 8'b00000000 ;
			15'h00001FCE : data <= 8'b00000000 ;
			15'h00001FCF : data <= 8'b00000000 ;
			15'h00001FD0 : data <= 8'b00000000 ;
			15'h00001FD1 : data <= 8'b00000000 ;
			15'h00001FD2 : data <= 8'b00000000 ;
			15'h00001FD3 : data <= 8'b00000000 ;
			15'h00001FD4 : data <= 8'b00000000 ;
			15'h00001FD5 : data <= 8'b00000000 ;
			15'h00001FD6 : data <= 8'b00000000 ;
			15'h00001FD7 : data <= 8'b00000000 ;
			15'h00001FD8 : data <= 8'b00000000 ;
			15'h00001FD9 : data <= 8'b00000000 ;
			15'h00001FDA : data <= 8'b00000000 ;
			15'h00001FDB : data <= 8'b00000000 ;
			15'h00001FDC : data <= 8'b00000000 ;
			15'h00001FDD : data <= 8'b00000000 ;
			15'h00001FDE : data <= 8'b00000000 ;
			15'h00001FDF : data <= 8'b00000000 ;
			15'h00001FE0 : data <= 8'b00000000 ;
			15'h00001FE1 : data <= 8'b00000000 ;
			15'h00001FE2 : data <= 8'b00000000 ;
			15'h00001FE3 : data <= 8'b00000000 ;
			15'h00001FE4 : data <= 8'b00000000 ;
			15'h00001FE5 : data <= 8'b00000000 ;
			15'h00001FE6 : data <= 8'b00000000 ;
			15'h00001FE7 : data <= 8'b00000000 ;
			15'h00001FE8 : data <= 8'b00000000 ;
			15'h00001FE9 : data <= 8'b00000000 ;
			15'h00001FEA : data <= 8'b00000000 ;
			15'h00001FEB : data <= 8'b00000000 ;
			15'h00001FEC : data <= 8'b00000000 ;
			15'h00001FED : data <= 8'b00000000 ;
			15'h00001FEE : data <= 8'b00000000 ;
			15'h00001FEF : data <= 8'b00000000 ;
			15'h00001FF0 : data <= 8'b00000000 ;
			15'h00001FF1 : data <= 8'b00000000 ;
			15'h00001FF2 : data <= 8'b00000000 ;
			15'h00001FF3 : data <= 8'b00000000 ;
			15'h00001FF4 : data <= 8'b00000000 ;
			15'h00001FF5 : data <= 8'b00000000 ;
			15'h00001FF6 : data <= 8'b00000000 ;
			15'h00001FF7 : data <= 8'b00000000 ;
			15'h00001FF8 : data <= 8'b00000000 ;
			15'h00001FF9 : data <= 8'b00000000 ;
			15'h00001FFA : data <= 8'b00000000 ;
			15'h00001FFB : data <= 8'b00000000 ;
			15'h00001FFC : data <= 8'b00000000 ;
			15'h00001FFD : data <= 8'b00000000 ;
			15'h00001FFE : data <= 8'b00000000 ;
			15'h00001FFF : data <= 8'b00000000 ;
			15'h00002000 : data <= 8'b00000000 ;
			15'h00002001 : data <= 8'b00000000 ;
			15'h00002002 : data <= 8'b00000000 ;
			15'h00002003 : data <= 8'b00000000 ;
			15'h00002004 : data <= 8'b00000000 ;
			15'h00002005 : data <= 8'b00000000 ;
			15'h00002006 : data <= 8'b00000000 ;
			15'h00002007 : data <= 8'b00000000 ;
			15'h00002008 : data <= 8'b00000000 ;
			15'h00002009 : data <= 8'b00000000 ;
			15'h0000200A : data <= 8'b00000000 ;
			15'h0000200B : data <= 8'b00000000 ;
			15'h0000200C : data <= 8'b00000000 ;
			15'h0000200D : data <= 8'b00000000 ;
			15'h0000200E : data <= 8'b00000000 ;
			15'h0000200F : data <= 8'b00000000 ;
			15'h00002010 : data <= 8'b00000000 ;
			15'h00002011 : data <= 8'b00000000 ;
			15'h00002012 : data <= 8'b00000000 ;
			15'h00002013 : data <= 8'b00000000 ;
			15'h00002014 : data <= 8'b00000000 ;
			15'h00002015 : data <= 8'b00000000 ;
			15'h00002016 : data <= 8'b00000000 ;
			15'h00002017 : data <= 8'b00000000 ;
			15'h00002018 : data <= 8'b00000000 ;
			15'h00002019 : data <= 8'b00000000 ;
			15'h0000201A : data <= 8'b00000000 ;
			15'h0000201B : data <= 8'b00000000 ;
			15'h0000201C : data <= 8'b00000000 ;
			15'h0000201D : data <= 8'b00000000 ;
			15'h0000201E : data <= 8'b00000000 ;
			15'h0000201F : data <= 8'b00000000 ;
			15'h00002020 : data <= 8'b00000000 ;
			15'h00002021 : data <= 8'b00000000 ;
			15'h00002022 : data <= 8'b00000000 ;
			15'h00002023 : data <= 8'b00000000 ;
			15'h00002024 : data <= 8'b00000000 ;
			15'h00002025 : data <= 8'b00000000 ;
			15'h00002026 : data <= 8'b00000000 ;
			15'h00002027 : data <= 8'b00000000 ;
			15'h00002028 : data <= 8'b00000000 ;
			15'h00002029 : data <= 8'b00000000 ;
			15'h0000202A : data <= 8'b00000000 ;
			15'h0000202B : data <= 8'b00000000 ;
			15'h0000202C : data <= 8'b00000000 ;
			15'h0000202D : data <= 8'b00000000 ;
			15'h0000202E : data <= 8'b00000000 ;
			15'h0000202F : data <= 8'b00000000 ;
			15'h00002030 : data <= 8'b00000000 ;
			15'h00002031 : data <= 8'b00000000 ;
			15'h00002032 : data <= 8'b00000000 ;
			15'h00002033 : data <= 8'b00000000 ;
			15'h00002034 : data <= 8'b00000000 ;
			15'h00002035 : data <= 8'b00000000 ;
			15'h00002036 : data <= 8'b00000000 ;
			15'h00002037 : data <= 8'b00000000 ;
			15'h00002038 : data <= 8'b00000000 ;
			15'h00002039 : data <= 8'b00000000 ;
			15'h0000203A : data <= 8'b00000000 ;
			15'h0000203B : data <= 8'b00000000 ;
			15'h0000203C : data <= 8'b00000000 ;
			15'h0000203D : data <= 8'b00000000 ;
			15'h0000203E : data <= 8'b00000000 ;
			15'h0000203F : data <= 8'b00000000 ;
			15'h00002040 : data <= 8'b00000000 ;
			15'h00002041 : data <= 8'b00000000 ;
			15'h00002042 : data <= 8'b00000000 ;
			15'h00002043 : data <= 8'b00000000 ;
			15'h00002044 : data <= 8'b00000000 ;
			15'h00002045 : data <= 8'b00000000 ;
			15'h00002046 : data <= 8'b00000000 ;
			15'h00002047 : data <= 8'b00000000 ;
			15'h00002048 : data <= 8'b00000000 ;
			15'h00002049 : data <= 8'b00000000 ;
			15'h0000204A : data <= 8'b00000000 ;
			15'h0000204B : data <= 8'b00000000 ;
			15'h0000204C : data <= 8'b00000000 ;
			15'h0000204D : data <= 8'b00000000 ;
			15'h0000204E : data <= 8'b00000000 ;
			15'h0000204F : data <= 8'b00000000 ;
			15'h00002050 : data <= 8'b00000000 ;
			15'h00002051 : data <= 8'b00000000 ;
			15'h00002052 : data <= 8'b00000000 ;
			15'h00002053 : data <= 8'b00000000 ;
			15'h00002054 : data <= 8'b00000000 ;
			15'h00002055 : data <= 8'b00000000 ;
			15'h00002056 : data <= 8'b00000000 ;
			15'h00002057 : data <= 8'b00000000 ;
			15'h00002058 : data <= 8'b00000000 ;
			15'h00002059 : data <= 8'b00000000 ;
			15'h0000205A : data <= 8'b00000000 ;
			15'h0000205B : data <= 8'b00000000 ;
			15'h0000205C : data <= 8'b00000000 ;
			15'h0000205D : data <= 8'b00000000 ;
			15'h0000205E : data <= 8'b00000000 ;
			15'h0000205F : data <= 8'b00000000 ;
			15'h00002060 : data <= 8'b00000000 ;
			15'h00002061 : data <= 8'b00000000 ;
			15'h00002062 : data <= 8'b00000000 ;
			15'h00002063 : data <= 8'b00000000 ;
			15'h00002064 : data <= 8'b00000000 ;
			15'h00002065 : data <= 8'b00000000 ;
			15'h00002066 : data <= 8'b00000000 ;
			15'h00002067 : data <= 8'b00000000 ;
			15'h00002068 : data <= 8'b00000000 ;
			15'h00002069 : data <= 8'b00000000 ;
			15'h0000206A : data <= 8'b00000000 ;
			15'h0000206B : data <= 8'b00000000 ;
			15'h0000206C : data <= 8'b00000000 ;
			15'h0000206D : data <= 8'b00000000 ;
			15'h0000206E : data <= 8'b00000000 ;
			15'h0000206F : data <= 8'b00000000 ;
			15'h00002070 : data <= 8'b00000000 ;
			15'h00002071 : data <= 8'b00000000 ;
			15'h00002072 : data <= 8'b00000000 ;
			15'h00002073 : data <= 8'b00000000 ;
			15'h00002074 : data <= 8'b00000000 ;
			15'h00002075 : data <= 8'b00000000 ;
			15'h00002076 : data <= 8'b00000000 ;
			15'h00002077 : data <= 8'b00000000 ;
			15'h00002078 : data <= 8'b00000000 ;
			15'h00002079 : data <= 8'b00000000 ;
			15'h0000207A : data <= 8'b00000000 ;
			15'h0000207B : data <= 8'b00000000 ;
			15'h0000207C : data <= 8'b00000000 ;
			15'h0000207D : data <= 8'b00000000 ;
			15'h0000207E : data <= 8'b00000000 ;
			15'h0000207F : data <= 8'b00000000 ;
			15'h00002080 : data <= 8'b00000000 ;
			15'h00002081 : data <= 8'b00000000 ;
			15'h00002082 : data <= 8'b00000000 ;
			15'h00002083 : data <= 8'b00000000 ;
			15'h00002084 : data <= 8'b00000000 ;
			15'h00002085 : data <= 8'b00000000 ;
			15'h00002086 : data <= 8'b00000000 ;
			15'h00002087 : data <= 8'b00000000 ;
			15'h00002088 : data <= 8'b00000000 ;
			15'h00002089 : data <= 8'b00000000 ;
			15'h0000208A : data <= 8'b00000000 ;
			15'h0000208B : data <= 8'b00000000 ;
			15'h0000208C : data <= 8'b00000000 ;
			15'h0000208D : data <= 8'b00000000 ;
			15'h0000208E : data <= 8'b00000000 ;
			15'h0000208F : data <= 8'b00000000 ;
			15'h00002090 : data <= 8'b00000000 ;
			15'h00002091 : data <= 8'b00000000 ;
			15'h00002092 : data <= 8'b00000000 ;
			15'h00002093 : data <= 8'b00000000 ;
			15'h00002094 : data <= 8'b00000000 ;
			15'h00002095 : data <= 8'b00000000 ;
			15'h00002096 : data <= 8'b00000000 ;
			15'h00002097 : data <= 8'b00000000 ;
			15'h00002098 : data <= 8'b00000000 ;
			15'h00002099 : data <= 8'b00000000 ;
			15'h0000209A : data <= 8'b00000000 ;
			15'h0000209B : data <= 8'b00000000 ;
			15'h0000209C : data <= 8'b00000000 ;
			15'h0000209D : data <= 8'b00000000 ;
			15'h0000209E : data <= 8'b00000000 ;
			15'h0000209F : data <= 8'b00000000 ;
			15'h000020A0 : data <= 8'b00000000 ;
			15'h000020A1 : data <= 8'b00000000 ;
			15'h000020A2 : data <= 8'b00000000 ;
			15'h000020A3 : data <= 8'b00000000 ;
			15'h000020A4 : data <= 8'b00000000 ;
			15'h000020A5 : data <= 8'b00000000 ;
			15'h000020A6 : data <= 8'b00000000 ;
			15'h000020A7 : data <= 8'b00000000 ;
			15'h000020A8 : data <= 8'b00000000 ;
			15'h000020A9 : data <= 8'b00000000 ;
			15'h000020AA : data <= 8'b00000000 ;
			15'h000020AB : data <= 8'b00000000 ;
			15'h000020AC : data <= 8'b00000000 ;
			15'h000020AD : data <= 8'b00000000 ;
			15'h000020AE : data <= 8'b00000000 ;
			15'h000020AF : data <= 8'b00000000 ;
			15'h000020B0 : data <= 8'b00000000 ;
			15'h000020B1 : data <= 8'b00000000 ;
			15'h000020B2 : data <= 8'b00000000 ;
			15'h000020B3 : data <= 8'b00000000 ;
			15'h000020B4 : data <= 8'b00000000 ;
			15'h000020B5 : data <= 8'b00000000 ;
			15'h000020B6 : data <= 8'b00000000 ;
			15'h000020B7 : data <= 8'b00000000 ;
			15'h000020B8 : data <= 8'b00000000 ;
			15'h000020B9 : data <= 8'b00000000 ;
			15'h000020BA : data <= 8'b00000000 ;
			15'h000020BB : data <= 8'b00000000 ;
			15'h000020BC : data <= 8'b00000000 ;
			15'h000020BD : data <= 8'b00000000 ;
			15'h000020BE : data <= 8'b00000000 ;
			15'h000020BF : data <= 8'b00000000 ;
			15'h000020C0 : data <= 8'b00000000 ;
			15'h000020C1 : data <= 8'b00000000 ;
			15'h000020C2 : data <= 8'b00000000 ;
			15'h000020C3 : data <= 8'b00000000 ;
			15'h000020C4 : data <= 8'b00000000 ;
			15'h000020C5 : data <= 8'b00000000 ;
			15'h000020C6 : data <= 8'b00000000 ;
			15'h000020C7 : data <= 8'b00000000 ;
			15'h000020C8 : data <= 8'b00000000 ;
			15'h000020C9 : data <= 8'b00000000 ;
			15'h000020CA : data <= 8'b00000000 ;
			15'h000020CB : data <= 8'b00000000 ;
			15'h000020CC : data <= 8'b00000000 ;
			15'h000020CD : data <= 8'b00000000 ;
			15'h000020CE : data <= 8'b00000000 ;
			15'h000020CF : data <= 8'b00000000 ;
			15'h000020D0 : data <= 8'b00000000 ;
			15'h000020D1 : data <= 8'b00000000 ;
			15'h000020D2 : data <= 8'b00000000 ;
			15'h000020D3 : data <= 8'b00000000 ;
			15'h000020D4 : data <= 8'b00000000 ;
			15'h000020D5 : data <= 8'b00000000 ;
			15'h000020D6 : data <= 8'b00000000 ;
			15'h000020D7 : data <= 8'b00000000 ;
			15'h000020D8 : data <= 8'b00000000 ;
			15'h000020D9 : data <= 8'b00000000 ;
			15'h000020DA : data <= 8'b00000000 ;
			15'h000020DB : data <= 8'b00000000 ;
			15'h000020DC : data <= 8'b00000000 ;
			15'h000020DD : data <= 8'b00000000 ;
			15'h000020DE : data <= 8'b00000000 ;
			15'h000020DF : data <= 8'b00000000 ;
			15'h000020E0 : data <= 8'b00000000 ;
			15'h000020E1 : data <= 8'b00000000 ;
			15'h000020E2 : data <= 8'b00000000 ;
			15'h000020E3 : data <= 8'b00000000 ;
			15'h000020E4 : data <= 8'b00000000 ;
			15'h000020E5 : data <= 8'b00000000 ;
			15'h000020E6 : data <= 8'b00000000 ;
			15'h000020E7 : data <= 8'b00000000 ;
			15'h000020E8 : data <= 8'b00000000 ;
			15'h000020E9 : data <= 8'b00000000 ;
			15'h000020EA : data <= 8'b00000000 ;
			15'h000020EB : data <= 8'b00000000 ;
			15'h000020EC : data <= 8'b00000000 ;
			15'h000020ED : data <= 8'b00000000 ;
			15'h000020EE : data <= 8'b00000000 ;
			15'h000020EF : data <= 8'b00000000 ;
			15'h000020F0 : data <= 8'b00000000 ;
			15'h000020F1 : data <= 8'b00000000 ;
			15'h000020F2 : data <= 8'b00000000 ;
			15'h000020F3 : data <= 8'b00000000 ;
			15'h000020F4 : data <= 8'b00000000 ;
			15'h000020F5 : data <= 8'b00000000 ;
			15'h000020F6 : data <= 8'b00000000 ;
			15'h000020F7 : data <= 8'b00000000 ;
			15'h000020F8 : data <= 8'b00000000 ;
			15'h000020F9 : data <= 8'b00000000 ;
			15'h000020FA : data <= 8'b00000000 ;
			15'h000020FB : data <= 8'b00000000 ;
			15'h000020FC : data <= 8'b00000000 ;
			15'h000020FD : data <= 8'b00000000 ;
			15'h000020FE : data <= 8'b00000000 ;
			15'h000020FF : data <= 8'b00000000 ;
			15'h00002100 : data <= 8'b00000000 ;
			15'h00002101 : data <= 8'b00000000 ;
			15'h00002102 : data <= 8'b00000000 ;
			15'h00002103 : data <= 8'b00000000 ;
			15'h00002104 : data <= 8'b00000000 ;
			15'h00002105 : data <= 8'b00000000 ;
			15'h00002106 : data <= 8'b00000000 ;
			15'h00002107 : data <= 8'b00000000 ;
			15'h00002108 : data <= 8'b00000000 ;
			15'h00002109 : data <= 8'b00000000 ;
			15'h0000210A : data <= 8'b00000000 ;
			15'h0000210B : data <= 8'b00000000 ;
			15'h0000210C : data <= 8'b00000000 ;
			15'h0000210D : data <= 8'b00000000 ;
			15'h0000210E : data <= 8'b00000000 ;
			15'h0000210F : data <= 8'b00000000 ;
			15'h00002110 : data <= 8'b00000000 ;
			15'h00002111 : data <= 8'b00000000 ;
			15'h00002112 : data <= 8'b00000000 ;
			15'h00002113 : data <= 8'b00000000 ;
			15'h00002114 : data <= 8'b00000000 ;
			15'h00002115 : data <= 8'b00000000 ;
			15'h00002116 : data <= 8'b00000000 ;
			15'h00002117 : data <= 8'b00000000 ;
			15'h00002118 : data <= 8'b00000000 ;
			15'h00002119 : data <= 8'b00000000 ;
			15'h0000211A : data <= 8'b00000000 ;
			15'h0000211B : data <= 8'b00000000 ;
			15'h0000211C : data <= 8'b00000000 ;
			15'h0000211D : data <= 8'b00000000 ;
			15'h0000211E : data <= 8'b00000000 ;
			15'h0000211F : data <= 8'b00000000 ;
			15'h00002120 : data <= 8'b00000000 ;
			15'h00002121 : data <= 8'b00000000 ;
			15'h00002122 : data <= 8'b00000000 ;
			15'h00002123 : data <= 8'b00000000 ;
			15'h00002124 : data <= 8'b00000000 ;
			15'h00002125 : data <= 8'b00000000 ;
			15'h00002126 : data <= 8'b00000000 ;
			15'h00002127 : data <= 8'b00000000 ;
			15'h00002128 : data <= 8'b00000000 ;
			15'h00002129 : data <= 8'b00000000 ;
			15'h0000212A : data <= 8'b00000000 ;
			15'h0000212B : data <= 8'b00000000 ;
			15'h0000212C : data <= 8'b00000000 ;
			15'h0000212D : data <= 8'b00000000 ;
			15'h0000212E : data <= 8'b00000000 ;
			15'h0000212F : data <= 8'b00000000 ;
			15'h00002130 : data <= 8'b00000000 ;
			15'h00002131 : data <= 8'b00000000 ;
			15'h00002132 : data <= 8'b00000000 ;
			15'h00002133 : data <= 8'b00000000 ;
			15'h00002134 : data <= 8'b00000000 ;
			15'h00002135 : data <= 8'b00000000 ;
			15'h00002136 : data <= 8'b00000000 ;
			15'h00002137 : data <= 8'b00000000 ;
			15'h00002138 : data <= 8'b00000000 ;
			15'h00002139 : data <= 8'b00000000 ;
			15'h0000213A : data <= 8'b00000000 ;
			15'h0000213B : data <= 8'b00000000 ;
			15'h0000213C : data <= 8'b00000000 ;
			15'h0000213D : data <= 8'b00000000 ;
			15'h0000213E : data <= 8'b00000000 ;
			15'h0000213F : data <= 8'b00000000 ;
			15'h00002140 : data <= 8'b00000000 ;
			15'h00002141 : data <= 8'b00000000 ;
			15'h00002142 : data <= 8'b00000000 ;
			15'h00002143 : data <= 8'b00000000 ;
			15'h00002144 : data <= 8'b00000000 ;
			15'h00002145 : data <= 8'b00000000 ;
			15'h00002146 : data <= 8'b00000000 ;
			15'h00002147 : data <= 8'b00000000 ;
			15'h00002148 : data <= 8'b00000000 ;
			15'h00002149 : data <= 8'b00000000 ;
			15'h0000214A : data <= 8'b00000000 ;
			15'h0000214B : data <= 8'b00000000 ;
			15'h0000214C : data <= 8'b00000000 ;
			15'h0000214D : data <= 8'b00000000 ;
			15'h0000214E : data <= 8'b00000000 ;
			15'h0000214F : data <= 8'b00000000 ;
			15'h00002150 : data <= 8'b00000000 ;
			15'h00002151 : data <= 8'b00000000 ;
			15'h00002152 : data <= 8'b00000000 ;
			15'h00002153 : data <= 8'b00000000 ;
			15'h00002154 : data <= 8'b00000000 ;
			15'h00002155 : data <= 8'b00000000 ;
			15'h00002156 : data <= 8'b00000000 ;
			15'h00002157 : data <= 8'b00000000 ;
			15'h00002158 : data <= 8'b00000000 ;
			15'h00002159 : data <= 8'b00000000 ;
			15'h0000215A : data <= 8'b00000000 ;
			15'h0000215B : data <= 8'b00000000 ;
			15'h0000215C : data <= 8'b00000000 ;
			15'h0000215D : data <= 8'b00000000 ;
			15'h0000215E : data <= 8'b00000000 ;
			15'h0000215F : data <= 8'b00000000 ;
			15'h00002160 : data <= 8'b00000000 ;
			15'h00002161 : data <= 8'b00000000 ;
			15'h00002162 : data <= 8'b00000000 ;
			15'h00002163 : data <= 8'b00000000 ;
			15'h00002164 : data <= 8'b00000000 ;
			15'h00002165 : data <= 8'b00000000 ;
			15'h00002166 : data <= 8'b00000000 ;
			15'h00002167 : data <= 8'b00000000 ;
			15'h00002168 : data <= 8'b00000000 ;
			15'h00002169 : data <= 8'b00000000 ;
			15'h0000216A : data <= 8'b00000000 ;
			15'h0000216B : data <= 8'b00000000 ;
			15'h0000216C : data <= 8'b00000000 ;
			15'h0000216D : data <= 8'b00000000 ;
			15'h0000216E : data <= 8'b00000000 ;
			15'h0000216F : data <= 8'b00000000 ;
			15'h00002170 : data <= 8'b00000000 ;
			15'h00002171 : data <= 8'b00000000 ;
			15'h00002172 : data <= 8'b00000000 ;
			15'h00002173 : data <= 8'b00000000 ;
			15'h00002174 : data <= 8'b00000000 ;
			15'h00002175 : data <= 8'b00000000 ;
			15'h00002176 : data <= 8'b00000000 ;
			15'h00002177 : data <= 8'b00000000 ;
			15'h00002178 : data <= 8'b00000000 ;
			15'h00002179 : data <= 8'b00000000 ;
			15'h0000217A : data <= 8'b00000000 ;
			15'h0000217B : data <= 8'b00000000 ;
			15'h0000217C : data <= 8'b00000000 ;
			15'h0000217D : data <= 8'b00000000 ;
			15'h0000217E : data <= 8'b00000000 ;
			15'h0000217F : data <= 8'b00000000 ;
			15'h00002180 : data <= 8'b00000000 ;
			15'h00002181 : data <= 8'b00000000 ;
			15'h00002182 : data <= 8'b00000000 ;
			15'h00002183 : data <= 8'b00000000 ;
			15'h00002184 : data <= 8'b00000000 ;
			15'h00002185 : data <= 8'b00000000 ;
			15'h00002186 : data <= 8'b00000000 ;
			15'h00002187 : data <= 8'b00000000 ;
			15'h00002188 : data <= 8'b00000000 ;
			15'h00002189 : data <= 8'b00000000 ;
			15'h0000218A : data <= 8'b00000000 ;
			15'h0000218B : data <= 8'b00000000 ;
			15'h0000218C : data <= 8'b00000000 ;
			15'h0000218D : data <= 8'b00000000 ;
			15'h0000218E : data <= 8'b00000000 ;
			15'h0000218F : data <= 8'b00000000 ;
			15'h00002190 : data <= 8'b00000000 ;
			15'h00002191 : data <= 8'b00000000 ;
			15'h00002192 : data <= 8'b00000000 ;
			15'h00002193 : data <= 8'b00000000 ;
			15'h00002194 : data <= 8'b00000000 ;
			15'h00002195 : data <= 8'b00000000 ;
			15'h00002196 : data <= 8'b00000000 ;
			15'h00002197 : data <= 8'b00000000 ;
			15'h00002198 : data <= 8'b00000000 ;
			15'h00002199 : data <= 8'b00000000 ;
			15'h0000219A : data <= 8'b00000000 ;
			15'h0000219B : data <= 8'b00000000 ;
			15'h0000219C : data <= 8'b00000000 ;
			15'h0000219D : data <= 8'b00000000 ;
			15'h0000219E : data <= 8'b00000000 ;
			15'h0000219F : data <= 8'b00000000 ;
			15'h000021A0 : data <= 8'b00000000 ;
			15'h000021A1 : data <= 8'b00000000 ;
			15'h000021A2 : data <= 8'b00000000 ;
			15'h000021A3 : data <= 8'b00000000 ;
			15'h000021A4 : data <= 8'b00000000 ;
			15'h000021A5 : data <= 8'b00000000 ;
			15'h000021A6 : data <= 8'b00000000 ;
			15'h000021A7 : data <= 8'b00000000 ;
			15'h000021A8 : data <= 8'b00000000 ;
			15'h000021A9 : data <= 8'b00000000 ;
			15'h000021AA : data <= 8'b00000000 ;
			15'h000021AB : data <= 8'b00000000 ;
			15'h000021AC : data <= 8'b00000000 ;
			15'h000021AD : data <= 8'b00000000 ;
			15'h000021AE : data <= 8'b00000000 ;
			15'h000021AF : data <= 8'b00000000 ;
			15'h000021B0 : data <= 8'b00000000 ;
			15'h000021B1 : data <= 8'b00000000 ;
			15'h000021B2 : data <= 8'b00000000 ;
			15'h000021B3 : data <= 8'b00000000 ;
			15'h000021B4 : data <= 8'b00000000 ;
			15'h000021B5 : data <= 8'b00000000 ;
			15'h000021B6 : data <= 8'b00000000 ;
			15'h000021B7 : data <= 8'b00000000 ;
			15'h000021B8 : data <= 8'b00000000 ;
			15'h000021B9 : data <= 8'b00000000 ;
			15'h000021BA : data <= 8'b00000000 ;
			15'h000021BB : data <= 8'b00000000 ;
			15'h000021BC : data <= 8'b00000000 ;
			15'h000021BD : data <= 8'b00000000 ;
			15'h000021BE : data <= 8'b00000000 ;
			15'h000021BF : data <= 8'b00000000 ;
			15'h000021C0 : data <= 8'b00000000 ;
			15'h000021C1 : data <= 8'b00000000 ;
			15'h000021C2 : data <= 8'b00000000 ;
			15'h000021C3 : data <= 8'b00000000 ;
			15'h000021C4 : data <= 8'b00000000 ;
			15'h000021C5 : data <= 8'b00000000 ;
			15'h000021C6 : data <= 8'b00000000 ;
			15'h000021C7 : data <= 8'b00000000 ;
			15'h000021C8 : data <= 8'b00000000 ;
			15'h000021C9 : data <= 8'b00000000 ;
			15'h000021CA : data <= 8'b00000000 ;
			15'h000021CB : data <= 8'b00000000 ;
			15'h000021CC : data <= 8'b00000000 ;
			15'h000021CD : data <= 8'b00000000 ;
			15'h000021CE : data <= 8'b00000000 ;
			15'h000021CF : data <= 8'b00000000 ;
			15'h000021D0 : data <= 8'b00000000 ;
			15'h000021D1 : data <= 8'b00000000 ;
			15'h000021D2 : data <= 8'b00000000 ;
			15'h000021D3 : data <= 8'b00000000 ;
			15'h000021D4 : data <= 8'b00000000 ;
			15'h000021D5 : data <= 8'b00000000 ;
			15'h000021D6 : data <= 8'b00000000 ;
			15'h000021D7 : data <= 8'b00000000 ;
			15'h000021D8 : data <= 8'b00000000 ;
			15'h000021D9 : data <= 8'b00000000 ;
			15'h000021DA : data <= 8'b00000000 ;
			15'h000021DB : data <= 8'b00000000 ;
			15'h000021DC : data <= 8'b00000000 ;
			15'h000021DD : data <= 8'b00000000 ;
			15'h000021DE : data <= 8'b00000000 ;
			15'h000021DF : data <= 8'b00000000 ;
			15'h000021E0 : data <= 8'b00000000 ;
			15'h000021E1 : data <= 8'b00000000 ;
			15'h000021E2 : data <= 8'b00000000 ;
			15'h000021E3 : data <= 8'b00000000 ;
			15'h000021E4 : data <= 8'b00000000 ;
			15'h000021E5 : data <= 8'b00000000 ;
			15'h000021E6 : data <= 8'b00000000 ;
			15'h000021E7 : data <= 8'b00000000 ;
			15'h000021E8 : data <= 8'b00000000 ;
			15'h000021E9 : data <= 8'b00000000 ;
			15'h000021EA : data <= 8'b00000000 ;
			15'h000021EB : data <= 8'b00000000 ;
			15'h000021EC : data <= 8'b00000000 ;
			15'h000021ED : data <= 8'b00000000 ;
			15'h000021EE : data <= 8'b00000000 ;
			15'h000021EF : data <= 8'b00000000 ;
			15'h000021F0 : data <= 8'b00000000 ;
			15'h000021F1 : data <= 8'b00000000 ;
			15'h000021F2 : data <= 8'b00000000 ;
			15'h000021F3 : data <= 8'b00000000 ;
			15'h000021F4 : data <= 8'b00000000 ;
			15'h000021F5 : data <= 8'b00000000 ;
			15'h000021F6 : data <= 8'b00000000 ;
			15'h000021F7 : data <= 8'b00000000 ;
			15'h000021F8 : data <= 8'b00000000 ;
			15'h000021F9 : data <= 8'b00000000 ;
			15'h000021FA : data <= 8'b00000000 ;
			15'h000021FB : data <= 8'b00000000 ;
			15'h000021FC : data <= 8'b00000000 ;
			15'h000021FD : data <= 8'b00000000 ;
			15'h000021FE : data <= 8'b00000000 ;
			15'h000021FF : data <= 8'b00000000 ;
			15'h00002200 : data <= 8'b00000000 ;
			15'h00002201 : data <= 8'b00000000 ;
			15'h00002202 : data <= 8'b00000000 ;
			15'h00002203 : data <= 8'b00000000 ;
			15'h00002204 : data <= 8'b00000000 ;
			15'h00002205 : data <= 8'b00000000 ;
			15'h00002206 : data <= 8'b00000000 ;
			15'h00002207 : data <= 8'b00000000 ;
			15'h00002208 : data <= 8'b00000000 ;
			15'h00002209 : data <= 8'b00000000 ;
			15'h0000220A : data <= 8'b00000000 ;
			15'h0000220B : data <= 8'b00000000 ;
			15'h0000220C : data <= 8'b00000000 ;
			15'h0000220D : data <= 8'b00000000 ;
			15'h0000220E : data <= 8'b00000000 ;
			15'h0000220F : data <= 8'b00000000 ;
			15'h00002210 : data <= 8'b00000000 ;
			15'h00002211 : data <= 8'b00000000 ;
			15'h00002212 : data <= 8'b00000000 ;
			15'h00002213 : data <= 8'b00000000 ;
			15'h00002214 : data <= 8'b00000000 ;
			15'h00002215 : data <= 8'b00000000 ;
			15'h00002216 : data <= 8'b00000000 ;
			15'h00002217 : data <= 8'b00000000 ;
			15'h00002218 : data <= 8'b00000000 ;
			15'h00002219 : data <= 8'b00000000 ;
			15'h0000221A : data <= 8'b00000000 ;
			15'h0000221B : data <= 8'b00000000 ;
			15'h0000221C : data <= 8'b00000000 ;
			15'h0000221D : data <= 8'b00000000 ;
			15'h0000221E : data <= 8'b00000000 ;
			15'h0000221F : data <= 8'b00000000 ;
			15'h00002220 : data <= 8'b00000000 ;
			15'h00002221 : data <= 8'b00000000 ;
			15'h00002222 : data <= 8'b00000000 ;
			15'h00002223 : data <= 8'b00000000 ;
			15'h00002224 : data <= 8'b00000000 ;
			15'h00002225 : data <= 8'b00000000 ;
			15'h00002226 : data <= 8'b00000000 ;
			15'h00002227 : data <= 8'b00000000 ;
			15'h00002228 : data <= 8'b00000000 ;
			15'h00002229 : data <= 8'b00000000 ;
			15'h0000222A : data <= 8'b00000000 ;
			15'h0000222B : data <= 8'b00000000 ;
			15'h0000222C : data <= 8'b00000000 ;
			15'h0000222D : data <= 8'b00000000 ;
			15'h0000222E : data <= 8'b00000000 ;
			15'h0000222F : data <= 8'b00000000 ;
			15'h00002230 : data <= 8'b00000000 ;
			15'h00002231 : data <= 8'b00000000 ;
			15'h00002232 : data <= 8'b00000000 ;
			15'h00002233 : data <= 8'b00000000 ;
			15'h00002234 : data <= 8'b00000000 ;
			15'h00002235 : data <= 8'b00000000 ;
			15'h00002236 : data <= 8'b00000000 ;
			15'h00002237 : data <= 8'b00000000 ;
			15'h00002238 : data <= 8'b00000000 ;
			15'h00002239 : data <= 8'b00000000 ;
			15'h0000223A : data <= 8'b00000000 ;
			15'h0000223B : data <= 8'b00000000 ;
			15'h0000223C : data <= 8'b00000000 ;
			15'h0000223D : data <= 8'b00000000 ;
			15'h0000223E : data <= 8'b00000000 ;
			15'h0000223F : data <= 8'b00000000 ;
			15'h00002240 : data <= 8'b00000000 ;
			15'h00002241 : data <= 8'b00000000 ;
			15'h00002242 : data <= 8'b00000000 ;
			15'h00002243 : data <= 8'b00000000 ;
			15'h00002244 : data <= 8'b00000000 ;
			15'h00002245 : data <= 8'b00000000 ;
			15'h00002246 : data <= 8'b00000000 ;
			15'h00002247 : data <= 8'b00000000 ;
			15'h00002248 : data <= 8'b00000000 ;
			15'h00002249 : data <= 8'b00000000 ;
			15'h0000224A : data <= 8'b00000000 ;
			15'h0000224B : data <= 8'b00000000 ;
			15'h0000224C : data <= 8'b00000000 ;
			15'h0000224D : data <= 8'b00000000 ;
			15'h0000224E : data <= 8'b00000000 ;
			15'h0000224F : data <= 8'b00000000 ;
			15'h00002250 : data <= 8'b00000000 ;
			15'h00002251 : data <= 8'b00000000 ;
			15'h00002252 : data <= 8'b00000000 ;
			15'h00002253 : data <= 8'b00000000 ;
			15'h00002254 : data <= 8'b00000000 ;
			15'h00002255 : data <= 8'b00000000 ;
			15'h00002256 : data <= 8'b00000000 ;
			15'h00002257 : data <= 8'b00000000 ;
			15'h00002258 : data <= 8'b00000000 ;
			15'h00002259 : data <= 8'b00000000 ;
			15'h0000225A : data <= 8'b00000000 ;
			15'h0000225B : data <= 8'b00000000 ;
			15'h0000225C : data <= 8'b00000000 ;
			15'h0000225D : data <= 8'b00000000 ;
			15'h0000225E : data <= 8'b00000000 ;
			15'h0000225F : data <= 8'b00000000 ;
			15'h00002260 : data <= 8'b00000000 ;
			15'h00002261 : data <= 8'b00000000 ;
			15'h00002262 : data <= 8'b00000000 ;
			15'h00002263 : data <= 8'b00000000 ;
			15'h00002264 : data <= 8'b00000000 ;
			15'h00002265 : data <= 8'b00000000 ;
			15'h00002266 : data <= 8'b00000000 ;
			15'h00002267 : data <= 8'b00000000 ;
			15'h00002268 : data <= 8'b00000000 ;
			15'h00002269 : data <= 8'b00000000 ;
			15'h0000226A : data <= 8'b00000000 ;
			15'h0000226B : data <= 8'b00000000 ;
			15'h0000226C : data <= 8'b00000000 ;
			15'h0000226D : data <= 8'b00000000 ;
			15'h0000226E : data <= 8'b00000000 ;
			15'h0000226F : data <= 8'b00000000 ;
			15'h00002270 : data <= 8'b00000000 ;
			15'h00002271 : data <= 8'b00000000 ;
			15'h00002272 : data <= 8'b00000000 ;
			15'h00002273 : data <= 8'b00000000 ;
			15'h00002274 : data <= 8'b00000000 ;
			15'h00002275 : data <= 8'b00000000 ;
			15'h00002276 : data <= 8'b00000000 ;
			15'h00002277 : data <= 8'b00000000 ;
			15'h00002278 : data <= 8'b00000000 ;
			15'h00002279 : data <= 8'b00000000 ;
			15'h0000227A : data <= 8'b00000000 ;
			15'h0000227B : data <= 8'b00000000 ;
			15'h0000227C : data <= 8'b00000000 ;
			15'h0000227D : data <= 8'b00000000 ;
			15'h0000227E : data <= 8'b00000000 ;
			15'h0000227F : data <= 8'b00000000 ;
			15'h00002280 : data <= 8'b00000000 ;
			15'h00002281 : data <= 8'b00000000 ;
			15'h00002282 : data <= 8'b00000000 ;
			15'h00002283 : data <= 8'b00000000 ;
			15'h00002284 : data <= 8'b00000000 ;
			15'h00002285 : data <= 8'b00000000 ;
			15'h00002286 : data <= 8'b00000000 ;
			15'h00002287 : data <= 8'b00000000 ;
			15'h00002288 : data <= 8'b00000000 ;
			15'h00002289 : data <= 8'b00000000 ;
			15'h0000228A : data <= 8'b00000000 ;
			15'h0000228B : data <= 8'b00000000 ;
			15'h0000228C : data <= 8'b00000000 ;
			15'h0000228D : data <= 8'b00000000 ;
			15'h0000228E : data <= 8'b00000000 ;
			15'h0000228F : data <= 8'b00000000 ;
			15'h00002290 : data <= 8'b00000000 ;
			15'h00002291 : data <= 8'b00000000 ;
			15'h00002292 : data <= 8'b00000000 ;
			15'h00002293 : data <= 8'b00000000 ;
			15'h00002294 : data <= 8'b00000000 ;
			15'h00002295 : data <= 8'b00000000 ;
			15'h00002296 : data <= 8'b00000000 ;
			15'h00002297 : data <= 8'b00000000 ;
			15'h00002298 : data <= 8'b00000000 ;
			15'h00002299 : data <= 8'b00000000 ;
			15'h0000229A : data <= 8'b00000000 ;
			15'h0000229B : data <= 8'b00000000 ;
			15'h0000229C : data <= 8'b00000000 ;
			15'h0000229D : data <= 8'b00000000 ;
			15'h0000229E : data <= 8'b00000000 ;
			15'h0000229F : data <= 8'b00000000 ;
			15'h000022A0 : data <= 8'b00000000 ;
			15'h000022A1 : data <= 8'b00000000 ;
			15'h000022A2 : data <= 8'b00000000 ;
			15'h000022A3 : data <= 8'b00000000 ;
			15'h000022A4 : data <= 8'b00000000 ;
			15'h000022A5 : data <= 8'b00000000 ;
			15'h000022A6 : data <= 8'b00000000 ;
			15'h000022A7 : data <= 8'b00000000 ;
			15'h000022A8 : data <= 8'b00000000 ;
			15'h000022A9 : data <= 8'b00000000 ;
			15'h000022AA : data <= 8'b00000000 ;
			15'h000022AB : data <= 8'b00000000 ;
			15'h000022AC : data <= 8'b00000000 ;
			15'h000022AD : data <= 8'b00000000 ;
			15'h000022AE : data <= 8'b00000000 ;
			15'h000022AF : data <= 8'b00000000 ;
			15'h000022B0 : data <= 8'b00000000 ;
			15'h000022B1 : data <= 8'b00000000 ;
			15'h000022B2 : data <= 8'b00000000 ;
			15'h000022B3 : data <= 8'b00000000 ;
			15'h000022B4 : data <= 8'b00000000 ;
			15'h000022B5 : data <= 8'b00000000 ;
			15'h000022B6 : data <= 8'b00000000 ;
			15'h000022B7 : data <= 8'b00000000 ;
			15'h000022B8 : data <= 8'b00000000 ;
			15'h000022B9 : data <= 8'b00000000 ;
			15'h000022BA : data <= 8'b00000000 ;
			15'h000022BB : data <= 8'b00000000 ;
			15'h000022BC : data <= 8'b00000000 ;
			15'h000022BD : data <= 8'b00000000 ;
			15'h000022BE : data <= 8'b00000000 ;
			15'h000022BF : data <= 8'b00000000 ;
			15'h000022C0 : data <= 8'b00000000 ;
			15'h000022C1 : data <= 8'b00000000 ;
			15'h000022C2 : data <= 8'b00000000 ;
			15'h000022C3 : data <= 8'b00000000 ;
			15'h000022C4 : data <= 8'b00000000 ;
			15'h000022C5 : data <= 8'b00000000 ;
			15'h000022C6 : data <= 8'b00000000 ;
			15'h000022C7 : data <= 8'b00000000 ;
			15'h000022C8 : data <= 8'b00000000 ;
			15'h000022C9 : data <= 8'b00000000 ;
			15'h000022CA : data <= 8'b00000000 ;
			15'h000022CB : data <= 8'b00000000 ;
			15'h000022CC : data <= 8'b00000000 ;
			15'h000022CD : data <= 8'b00000000 ;
			15'h000022CE : data <= 8'b00000000 ;
			15'h000022CF : data <= 8'b00000000 ;
			15'h000022D0 : data <= 8'b00000000 ;
			15'h000022D1 : data <= 8'b00000000 ;
			15'h000022D2 : data <= 8'b00000000 ;
			15'h000022D3 : data <= 8'b00000000 ;
			15'h000022D4 : data <= 8'b00000000 ;
			15'h000022D5 : data <= 8'b00000000 ;
			15'h000022D6 : data <= 8'b00000000 ;
			15'h000022D7 : data <= 8'b00000000 ;
			15'h000022D8 : data <= 8'b00000000 ;
			15'h000022D9 : data <= 8'b00000000 ;
			15'h000022DA : data <= 8'b00000000 ;
			15'h000022DB : data <= 8'b00000000 ;
			15'h000022DC : data <= 8'b00000000 ;
			15'h000022DD : data <= 8'b00000000 ;
			15'h000022DE : data <= 8'b00000000 ;
			15'h000022DF : data <= 8'b00000000 ;
			15'h000022E0 : data <= 8'b00000000 ;
			15'h000022E1 : data <= 8'b00000000 ;
			15'h000022E2 : data <= 8'b00000000 ;
			15'h000022E3 : data <= 8'b00000000 ;
			15'h000022E4 : data <= 8'b00000000 ;
			15'h000022E5 : data <= 8'b00000000 ;
			15'h000022E6 : data <= 8'b00000000 ;
			15'h000022E7 : data <= 8'b00000000 ;
			15'h000022E8 : data <= 8'b00000000 ;
			15'h000022E9 : data <= 8'b00000000 ;
			15'h000022EA : data <= 8'b00000000 ;
			15'h000022EB : data <= 8'b00000000 ;
			15'h000022EC : data <= 8'b00000000 ;
			15'h000022ED : data <= 8'b00000000 ;
			15'h000022EE : data <= 8'b00000000 ;
			15'h000022EF : data <= 8'b00000000 ;
			15'h000022F0 : data <= 8'b00000000 ;
			15'h000022F1 : data <= 8'b00000000 ;
			15'h000022F2 : data <= 8'b00000000 ;
			15'h000022F3 : data <= 8'b00000000 ;
			15'h000022F4 : data <= 8'b00000000 ;
			15'h000022F5 : data <= 8'b00000000 ;
			15'h000022F6 : data <= 8'b00000000 ;
			15'h000022F7 : data <= 8'b00000000 ;
			15'h000022F8 : data <= 8'b00000000 ;
			15'h000022F9 : data <= 8'b00000000 ;
			15'h000022FA : data <= 8'b00000000 ;
			15'h000022FB : data <= 8'b00000000 ;
			15'h000022FC : data <= 8'b00000000 ;
			15'h000022FD : data <= 8'b00000000 ;
			15'h000022FE : data <= 8'b00000000 ;
			15'h000022FF : data <= 8'b00000000 ;
			15'h00002300 : data <= 8'b00000000 ;
			15'h00002301 : data <= 8'b00000000 ;
			15'h00002302 : data <= 8'b00000000 ;
			15'h00002303 : data <= 8'b00000000 ;
			15'h00002304 : data <= 8'b00000000 ;
			15'h00002305 : data <= 8'b00000000 ;
			15'h00002306 : data <= 8'b00000000 ;
			15'h00002307 : data <= 8'b00000000 ;
			15'h00002308 : data <= 8'b00000000 ;
			15'h00002309 : data <= 8'b00000000 ;
			15'h0000230A : data <= 8'b00000000 ;
			15'h0000230B : data <= 8'b00000000 ;
			15'h0000230C : data <= 8'b00000000 ;
			15'h0000230D : data <= 8'b00000000 ;
			15'h0000230E : data <= 8'b00000000 ;
			15'h0000230F : data <= 8'b00000000 ;
			15'h00002310 : data <= 8'b00000000 ;
			15'h00002311 : data <= 8'b00000000 ;
			15'h00002312 : data <= 8'b00000000 ;
			15'h00002313 : data <= 8'b00000000 ;
			15'h00002314 : data <= 8'b00000000 ;
			15'h00002315 : data <= 8'b00000000 ;
			15'h00002316 : data <= 8'b00000000 ;
			15'h00002317 : data <= 8'b00000000 ;
			15'h00002318 : data <= 8'b00000000 ;
			15'h00002319 : data <= 8'b00000000 ;
			15'h0000231A : data <= 8'b00000000 ;
			15'h0000231B : data <= 8'b00000000 ;
			15'h0000231C : data <= 8'b00000000 ;
			15'h0000231D : data <= 8'b00000000 ;
			15'h0000231E : data <= 8'b00000000 ;
			15'h0000231F : data <= 8'b00000000 ;
			15'h00002320 : data <= 8'b00000000 ;
			15'h00002321 : data <= 8'b00000000 ;
			15'h00002322 : data <= 8'b00000000 ;
			15'h00002323 : data <= 8'b00000000 ;
			15'h00002324 : data <= 8'b00000000 ;
			15'h00002325 : data <= 8'b00000000 ;
			15'h00002326 : data <= 8'b00000000 ;
			15'h00002327 : data <= 8'b00000000 ;
			15'h00002328 : data <= 8'b00000000 ;
			15'h00002329 : data <= 8'b00000000 ;
			15'h0000232A : data <= 8'b00000000 ;
			15'h0000232B : data <= 8'b00000000 ;
			15'h0000232C : data <= 8'b00000000 ;
			15'h0000232D : data <= 8'b00000000 ;
			15'h0000232E : data <= 8'b00000000 ;
			15'h0000232F : data <= 8'b00000000 ;
			15'h00002330 : data <= 8'b00000000 ;
			15'h00002331 : data <= 8'b00000000 ;
			15'h00002332 : data <= 8'b00000000 ;
			15'h00002333 : data <= 8'b00000000 ;
			15'h00002334 : data <= 8'b00000000 ;
			15'h00002335 : data <= 8'b00000000 ;
			15'h00002336 : data <= 8'b00000000 ;
			15'h00002337 : data <= 8'b00000000 ;
			15'h00002338 : data <= 8'b00000000 ;
			15'h00002339 : data <= 8'b00000000 ;
			15'h0000233A : data <= 8'b00000000 ;
			15'h0000233B : data <= 8'b00000000 ;
			15'h0000233C : data <= 8'b00000000 ;
			15'h0000233D : data <= 8'b00000000 ;
			15'h0000233E : data <= 8'b00000000 ;
			15'h0000233F : data <= 8'b00000000 ;
			15'h00002340 : data <= 8'b00000000 ;
			15'h00002341 : data <= 8'b00000000 ;
			15'h00002342 : data <= 8'b00000000 ;
			15'h00002343 : data <= 8'b00000000 ;
			15'h00002344 : data <= 8'b00000000 ;
			15'h00002345 : data <= 8'b00000000 ;
			15'h00002346 : data <= 8'b00000000 ;
			15'h00002347 : data <= 8'b00000000 ;
			15'h00002348 : data <= 8'b00000000 ;
			15'h00002349 : data <= 8'b00000000 ;
			15'h0000234A : data <= 8'b00000000 ;
			15'h0000234B : data <= 8'b00000000 ;
			15'h0000234C : data <= 8'b00000000 ;
			15'h0000234D : data <= 8'b00000000 ;
			15'h0000234E : data <= 8'b00000000 ;
			15'h0000234F : data <= 8'b00000000 ;
			15'h00002350 : data <= 8'b00000000 ;
			15'h00002351 : data <= 8'b00000000 ;
			15'h00002352 : data <= 8'b00000000 ;
			15'h00002353 : data <= 8'b00000000 ;
			15'h00002354 : data <= 8'b00000000 ;
			15'h00002355 : data <= 8'b00000000 ;
			15'h00002356 : data <= 8'b00000000 ;
			15'h00002357 : data <= 8'b00000000 ;
			15'h00002358 : data <= 8'b00000000 ;
			15'h00002359 : data <= 8'b00000000 ;
			15'h0000235A : data <= 8'b00000000 ;
			15'h0000235B : data <= 8'b00000000 ;
			15'h0000235C : data <= 8'b00000000 ;
			15'h0000235D : data <= 8'b00000000 ;
			15'h0000235E : data <= 8'b00000000 ;
			15'h0000235F : data <= 8'b00000000 ;
			15'h00002360 : data <= 8'b00000000 ;
			15'h00002361 : data <= 8'b00000000 ;
			15'h00002362 : data <= 8'b00000000 ;
			15'h00002363 : data <= 8'b00000000 ;
			15'h00002364 : data <= 8'b00000000 ;
			15'h00002365 : data <= 8'b00000000 ;
			15'h00002366 : data <= 8'b00000000 ;
			15'h00002367 : data <= 8'b00000000 ;
			15'h00002368 : data <= 8'b00000000 ;
			15'h00002369 : data <= 8'b00000000 ;
			15'h0000236A : data <= 8'b00000000 ;
			15'h0000236B : data <= 8'b00000000 ;
			15'h0000236C : data <= 8'b00000000 ;
			15'h0000236D : data <= 8'b00000000 ;
			15'h0000236E : data <= 8'b00000000 ;
			15'h0000236F : data <= 8'b00000000 ;
			15'h00002370 : data <= 8'b00000000 ;
			15'h00002371 : data <= 8'b00000000 ;
			15'h00002372 : data <= 8'b00000000 ;
			15'h00002373 : data <= 8'b00000000 ;
			15'h00002374 : data <= 8'b00000000 ;
			15'h00002375 : data <= 8'b00000000 ;
			15'h00002376 : data <= 8'b00000000 ;
			15'h00002377 : data <= 8'b00000000 ;
			15'h00002378 : data <= 8'b00000000 ;
			15'h00002379 : data <= 8'b00000000 ;
			15'h0000237A : data <= 8'b00000000 ;
			15'h0000237B : data <= 8'b00000000 ;
			15'h0000237C : data <= 8'b00000000 ;
			15'h0000237D : data <= 8'b00000000 ;
			15'h0000237E : data <= 8'b00000000 ;
			15'h0000237F : data <= 8'b00000000 ;
			15'h00002380 : data <= 8'b00000000 ;
			15'h00002381 : data <= 8'b00000000 ;
			15'h00002382 : data <= 8'b00000000 ;
			15'h00002383 : data <= 8'b00000000 ;
			15'h00002384 : data <= 8'b00000000 ;
			15'h00002385 : data <= 8'b00000000 ;
			15'h00002386 : data <= 8'b00000000 ;
			15'h00002387 : data <= 8'b00000000 ;
			15'h00002388 : data <= 8'b00000000 ;
			15'h00002389 : data <= 8'b00000000 ;
			15'h0000238A : data <= 8'b00000000 ;
			15'h0000238B : data <= 8'b00000000 ;
			15'h0000238C : data <= 8'b00000000 ;
			15'h0000238D : data <= 8'b00000000 ;
			15'h0000238E : data <= 8'b00000000 ;
			15'h0000238F : data <= 8'b00000000 ;
			15'h00002390 : data <= 8'b00000000 ;
			15'h00002391 : data <= 8'b00000000 ;
			15'h00002392 : data <= 8'b00000000 ;
			15'h00002393 : data <= 8'b00000000 ;
			15'h00002394 : data <= 8'b00000000 ;
			15'h00002395 : data <= 8'b00000000 ;
			15'h00002396 : data <= 8'b00000000 ;
			15'h00002397 : data <= 8'b00000000 ;
			15'h00002398 : data <= 8'b00000000 ;
			15'h00002399 : data <= 8'b00000000 ;
			15'h0000239A : data <= 8'b00000000 ;
			15'h0000239B : data <= 8'b00000000 ;
			15'h0000239C : data <= 8'b00000000 ;
			15'h0000239D : data <= 8'b00000000 ;
			15'h0000239E : data <= 8'b00000000 ;
			15'h0000239F : data <= 8'b00000000 ;
			15'h000023A0 : data <= 8'b00000000 ;
			15'h000023A1 : data <= 8'b00000000 ;
			15'h000023A2 : data <= 8'b00000000 ;
			15'h000023A3 : data <= 8'b00000000 ;
			15'h000023A4 : data <= 8'b00000000 ;
			15'h000023A5 : data <= 8'b00000000 ;
			15'h000023A6 : data <= 8'b00000000 ;
			15'h000023A7 : data <= 8'b00000000 ;
			15'h000023A8 : data <= 8'b00000000 ;
			15'h000023A9 : data <= 8'b00000000 ;
			15'h000023AA : data <= 8'b00000000 ;
			15'h000023AB : data <= 8'b00000000 ;
			15'h000023AC : data <= 8'b00000000 ;
			15'h000023AD : data <= 8'b00000000 ;
			15'h000023AE : data <= 8'b00000000 ;
			15'h000023AF : data <= 8'b00000000 ;
			15'h000023B0 : data <= 8'b00000000 ;
			15'h000023B1 : data <= 8'b00000000 ;
			15'h000023B2 : data <= 8'b00000000 ;
			15'h000023B3 : data <= 8'b00000000 ;
			15'h000023B4 : data <= 8'b00000000 ;
			15'h000023B5 : data <= 8'b00000000 ;
			15'h000023B6 : data <= 8'b00000000 ;
			15'h000023B7 : data <= 8'b00000000 ;
			15'h000023B8 : data <= 8'b00000000 ;
			15'h000023B9 : data <= 8'b00000000 ;
			15'h000023BA : data <= 8'b00000000 ;
			15'h000023BB : data <= 8'b00000000 ;
			15'h000023BC : data <= 8'b00000000 ;
			15'h000023BD : data <= 8'b00000000 ;
			15'h000023BE : data <= 8'b00000000 ;
			15'h000023BF : data <= 8'b00000000 ;
			15'h000023C0 : data <= 8'b00000000 ;
			15'h000023C1 : data <= 8'b00000000 ;
			15'h000023C2 : data <= 8'b00000000 ;
			15'h000023C3 : data <= 8'b00000000 ;
			15'h000023C4 : data <= 8'b00000000 ;
			15'h000023C5 : data <= 8'b00000000 ;
			15'h000023C6 : data <= 8'b00000000 ;
			15'h000023C7 : data <= 8'b00000000 ;
			15'h000023C8 : data <= 8'b00000000 ;
			15'h000023C9 : data <= 8'b00000000 ;
			15'h000023CA : data <= 8'b00000000 ;
			15'h000023CB : data <= 8'b00000000 ;
			15'h000023CC : data <= 8'b00000000 ;
			15'h000023CD : data <= 8'b00000000 ;
			15'h000023CE : data <= 8'b00000000 ;
			15'h000023CF : data <= 8'b00000000 ;
			15'h000023D0 : data <= 8'b00000000 ;
			15'h000023D1 : data <= 8'b00000000 ;
			15'h000023D2 : data <= 8'b00000000 ;
			15'h000023D3 : data <= 8'b00000000 ;
			15'h000023D4 : data <= 8'b00000000 ;
			15'h000023D5 : data <= 8'b00000000 ;
			15'h000023D6 : data <= 8'b00000000 ;
			15'h000023D7 : data <= 8'b00000000 ;
			15'h000023D8 : data <= 8'b00000000 ;
			15'h000023D9 : data <= 8'b00000000 ;
			15'h000023DA : data <= 8'b00000000 ;
			15'h000023DB : data <= 8'b00000000 ;
			15'h000023DC : data <= 8'b00000000 ;
			15'h000023DD : data <= 8'b00000000 ;
			15'h000023DE : data <= 8'b00000000 ;
			15'h000023DF : data <= 8'b00000000 ;
			15'h000023E0 : data <= 8'b00000000 ;
			15'h000023E1 : data <= 8'b00000000 ;
			15'h000023E2 : data <= 8'b00000000 ;
			15'h000023E3 : data <= 8'b00000000 ;
			15'h000023E4 : data <= 8'b00000000 ;
			15'h000023E5 : data <= 8'b00000000 ;
			15'h000023E6 : data <= 8'b00000000 ;
			15'h000023E7 : data <= 8'b00000000 ;
			15'h000023E8 : data <= 8'b00000000 ;
			15'h000023E9 : data <= 8'b00000000 ;
			15'h000023EA : data <= 8'b00000000 ;
			15'h000023EB : data <= 8'b00000000 ;
			15'h000023EC : data <= 8'b00000000 ;
			15'h000023ED : data <= 8'b00000000 ;
			15'h000023EE : data <= 8'b00000000 ;
			15'h000023EF : data <= 8'b00000000 ;
			15'h000023F0 : data <= 8'b00000000 ;
			15'h000023F1 : data <= 8'b00000000 ;
			15'h000023F2 : data <= 8'b00000000 ;
			15'h000023F3 : data <= 8'b00000000 ;
			15'h000023F4 : data <= 8'b00000000 ;
			15'h000023F5 : data <= 8'b00000000 ;
			15'h000023F6 : data <= 8'b00000000 ;
			15'h000023F7 : data <= 8'b00000000 ;
			15'h000023F8 : data <= 8'b00000000 ;
			15'h000023F9 : data <= 8'b00000000 ;
			15'h000023FA : data <= 8'b00000000 ;
			15'h000023FB : data <= 8'b00000000 ;
			15'h000023FC : data <= 8'b00000000 ;
			15'h000023FD : data <= 8'b00000000 ;
			15'h000023FE : data <= 8'b00000000 ;
			15'h000023FF : data <= 8'b00000000 ;
			15'h00002400 : data <= 8'b00000000 ;
			15'h00002401 : data <= 8'b00000000 ;
			15'h00002402 : data <= 8'b00000000 ;
			15'h00002403 : data <= 8'b00000000 ;
			15'h00002404 : data <= 8'b00000000 ;
			15'h00002405 : data <= 8'b00000000 ;
			15'h00002406 : data <= 8'b00000000 ;
			15'h00002407 : data <= 8'b00000000 ;
			15'h00002408 : data <= 8'b00000000 ;
			15'h00002409 : data <= 8'b00000000 ;
			15'h0000240A : data <= 8'b00000000 ;
			15'h0000240B : data <= 8'b00000000 ;
			15'h0000240C : data <= 8'b00000000 ;
			15'h0000240D : data <= 8'b00000000 ;
			15'h0000240E : data <= 8'b00000000 ;
			15'h0000240F : data <= 8'b00000000 ;
			15'h00002410 : data <= 8'b00000000 ;
			15'h00002411 : data <= 8'b00000000 ;
			15'h00002412 : data <= 8'b00000000 ;
			15'h00002413 : data <= 8'b00000000 ;
			15'h00002414 : data <= 8'b00000000 ;
			15'h00002415 : data <= 8'b00000000 ;
			15'h00002416 : data <= 8'b00000000 ;
			15'h00002417 : data <= 8'b00000000 ;
			15'h00002418 : data <= 8'b00000000 ;
			15'h00002419 : data <= 8'b00000000 ;
			15'h0000241A : data <= 8'b00000000 ;
			15'h0000241B : data <= 8'b00000000 ;
			15'h0000241C : data <= 8'b00000000 ;
			15'h0000241D : data <= 8'b00000000 ;
			15'h0000241E : data <= 8'b00000000 ;
			15'h0000241F : data <= 8'b00000000 ;
			15'h00002420 : data <= 8'b00000000 ;
			15'h00002421 : data <= 8'b00000000 ;
			15'h00002422 : data <= 8'b00000000 ;
			15'h00002423 : data <= 8'b00000000 ;
			15'h00002424 : data <= 8'b00000000 ;
			15'h00002425 : data <= 8'b00000000 ;
			15'h00002426 : data <= 8'b00000000 ;
			15'h00002427 : data <= 8'b00000000 ;
			15'h00002428 : data <= 8'b00000000 ;
			15'h00002429 : data <= 8'b00000000 ;
			15'h0000242A : data <= 8'b00000000 ;
			15'h0000242B : data <= 8'b00000000 ;
			15'h0000242C : data <= 8'b00000000 ;
			15'h0000242D : data <= 8'b00000000 ;
			15'h0000242E : data <= 8'b00000000 ;
			15'h0000242F : data <= 8'b00000000 ;
			15'h00002430 : data <= 8'b00000000 ;
			15'h00002431 : data <= 8'b00000000 ;
			15'h00002432 : data <= 8'b00000000 ;
			15'h00002433 : data <= 8'b00000000 ;
			15'h00002434 : data <= 8'b00000000 ;
			15'h00002435 : data <= 8'b00000000 ;
			15'h00002436 : data <= 8'b00000000 ;
			15'h00002437 : data <= 8'b00000000 ;
			15'h00002438 : data <= 8'b00000000 ;
			15'h00002439 : data <= 8'b00000000 ;
			15'h0000243A : data <= 8'b00000000 ;
			15'h0000243B : data <= 8'b00000000 ;
			15'h0000243C : data <= 8'b00000000 ;
			15'h0000243D : data <= 8'b00000000 ;
			15'h0000243E : data <= 8'b00000000 ;
			15'h0000243F : data <= 8'b00000000 ;
			15'h00002440 : data <= 8'b00000000 ;
			15'h00002441 : data <= 8'b00000000 ;
			15'h00002442 : data <= 8'b00000000 ;
			15'h00002443 : data <= 8'b00000000 ;
			15'h00002444 : data <= 8'b00000000 ;
			15'h00002445 : data <= 8'b00000000 ;
			15'h00002446 : data <= 8'b00000000 ;
			15'h00002447 : data <= 8'b00000000 ;
			15'h00002448 : data <= 8'b00000000 ;
			15'h00002449 : data <= 8'b00000000 ;
			15'h0000244A : data <= 8'b00000000 ;
			15'h0000244B : data <= 8'b00000000 ;
			15'h0000244C : data <= 8'b00000000 ;
			15'h0000244D : data <= 8'b00000000 ;
			15'h0000244E : data <= 8'b00000000 ;
			15'h0000244F : data <= 8'b00000000 ;
			15'h00002450 : data <= 8'b00000000 ;
			15'h00002451 : data <= 8'b00000000 ;
			15'h00002452 : data <= 8'b00000000 ;
			15'h00002453 : data <= 8'b00000000 ;
			15'h00002454 : data <= 8'b00000000 ;
			15'h00002455 : data <= 8'b00000000 ;
			15'h00002456 : data <= 8'b00000000 ;
			15'h00002457 : data <= 8'b00000000 ;
			15'h00002458 : data <= 8'b00000000 ;
			15'h00002459 : data <= 8'b00000000 ;
			15'h0000245A : data <= 8'b00000000 ;
			15'h0000245B : data <= 8'b00000000 ;
			15'h0000245C : data <= 8'b00000000 ;
			15'h0000245D : data <= 8'b00000000 ;
			15'h0000245E : data <= 8'b00000000 ;
			15'h0000245F : data <= 8'b00000000 ;
			15'h00002460 : data <= 8'b00000000 ;
			15'h00002461 : data <= 8'b00000000 ;
			15'h00002462 : data <= 8'b00000000 ;
			15'h00002463 : data <= 8'b00000000 ;
			15'h00002464 : data <= 8'b00000000 ;
			15'h00002465 : data <= 8'b00000000 ;
			15'h00002466 : data <= 8'b00000000 ;
			15'h00002467 : data <= 8'b00000000 ;
			15'h00002468 : data <= 8'b00000000 ;
			15'h00002469 : data <= 8'b00000000 ;
			15'h0000246A : data <= 8'b00000000 ;
			15'h0000246B : data <= 8'b00000000 ;
			15'h0000246C : data <= 8'b00000000 ;
			15'h0000246D : data <= 8'b00000000 ;
			15'h0000246E : data <= 8'b00000000 ;
			15'h0000246F : data <= 8'b00000000 ;
			15'h00002470 : data <= 8'b00000000 ;
			15'h00002471 : data <= 8'b00000000 ;
			15'h00002472 : data <= 8'b00000000 ;
			15'h00002473 : data <= 8'b00000000 ;
			15'h00002474 : data <= 8'b00000000 ;
			15'h00002475 : data <= 8'b00000000 ;
			15'h00002476 : data <= 8'b00000000 ;
			15'h00002477 : data <= 8'b00000000 ;
			15'h00002478 : data <= 8'b00000000 ;
			15'h00002479 : data <= 8'b00000000 ;
			15'h0000247A : data <= 8'b00000000 ;
			15'h0000247B : data <= 8'b00000000 ;
			15'h0000247C : data <= 8'b00000000 ;
			15'h0000247D : data <= 8'b00000000 ;
			15'h0000247E : data <= 8'b00000000 ;
			15'h0000247F : data <= 8'b00000000 ;
			15'h00002480 : data <= 8'b00000000 ;
			15'h00002481 : data <= 8'b00000000 ;
			15'h00002482 : data <= 8'b00000000 ;
			15'h00002483 : data <= 8'b00000000 ;
			15'h00002484 : data <= 8'b00000000 ;
			15'h00002485 : data <= 8'b00000000 ;
			15'h00002486 : data <= 8'b00000000 ;
			15'h00002487 : data <= 8'b00000000 ;
			15'h00002488 : data <= 8'b00000000 ;
			15'h00002489 : data <= 8'b00000000 ;
			15'h0000248A : data <= 8'b00000000 ;
			15'h0000248B : data <= 8'b00000000 ;
			15'h0000248C : data <= 8'b00000000 ;
			15'h0000248D : data <= 8'b00000000 ;
			15'h0000248E : data <= 8'b00000000 ;
			15'h0000248F : data <= 8'b00000000 ;
			15'h00002490 : data <= 8'b00000000 ;
			15'h00002491 : data <= 8'b00000000 ;
			15'h00002492 : data <= 8'b00000000 ;
			15'h00002493 : data <= 8'b00000000 ;
			15'h00002494 : data <= 8'b00000000 ;
			15'h00002495 : data <= 8'b00000000 ;
			15'h00002496 : data <= 8'b00000000 ;
			15'h00002497 : data <= 8'b00000000 ;
			15'h00002498 : data <= 8'b00000000 ;
			15'h00002499 : data <= 8'b00000000 ;
			15'h0000249A : data <= 8'b00000000 ;
			15'h0000249B : data <= 8'b00000000 ;
			15'h0000249C : data <= 8'b00000000 ;
			15'h0000249D : data <= 8'b00000000 ;
			15'h0000249E : data <= 8'b00000000 ;
			15'h0000249F : data <= 8'b00000000 ;
			15'h000024A0 : data <= 8'b00000000 ;
			15'h000024A1 : data <= 8'b00000000 ;
			15'h000024A2 : data <= 8'b00000000 ;
			15'h000024A3 : data <= 8'b00000000 ;
			15'h000024A4 : data <= 8'b00000000 ;
			15'h000024A5 : data <= 8'b00000000 ;
			15'h000024A6 : data <= 8'b00000000 ;
			15'h000024A7 : data <= 8'b00000000 ;
			15'h000024A8 : data <= 8'b00000000 ;
			15'h000024A9 : data <= 8'b00000000 ;
			15'h000024AA : data <= 8'b00000000 ;
			15'h000024AB : data <= 8'b00000000 ;
			15'h000024AC : data <= 8'b00000000 ;
			15'h000024AD : data <= 8'b00000000 ;
			15'h000024AE : data <= 8'b00000000 ;
			15'h000024AF : data <= 8'b00000000 ;
			15'h000024B0 : data <= 8'b00000000 ;
			15'h000024B1 : data <= 8'b00000000 ;
			15'h000024B2 : data <= 8'b00000000 ;
			15'h000024B3 : data <= 8'b00000000 ;
			15'h000024B4 : data <= 8'b00000000 ;
			15'h000024B5 : data <= 8'b00000000 ;
			15'h000024B6 : data <= 8'b00000000 ;
			15'h000024B7 : data <= 8'b00000000 ;
			15'h000024B8 : data <= 8'b00000000 ;
			15'h000024B9 : data <= 8'b00000000 ;
			15'h000024BA : data <= 8'b00000000 ;
			15'h000024BB : data <= 8'b00000000 ;
			15'h000024BC : data <= 8'b00000000 ;
			15'h000024BD : data <= 8'b00000000 ;
			15'h000024BE : data <= 8'b00000000 ;
			15'h000024BF : data <= 8'b00000000 ;
			15'h000024C0 : data <= 8'b00000000 ;
			15'h000024C1 : data <= 8'b00000000 ;
			15'h000024C2 : data <= 8'b00000000 ;
			15'h000024C3 : data <= 8'b00000000 ;
			15'h000024C4 : data <= 8'b00000000 ;
			15'h000024C5 : data <= 8'b00000000 ;
			15'h000024C6 : data <= 8'b00000000 ;
			15'h000024C7 : data <= 8'b00000000 ;
			15'h000024C8 : data <= 8'b00000000 ;
			15'h000024C9 : data <= 8'b00000000 ;
			15'h000024CA : data <= 8'b00000000 ;
			15'h000024CB : data <= 8'b00000000 ;
			15'h000024CC : data <= 8'b00000000 ;
			15'h000024CD : data <= 8'b00000000 ;
			15'h000024CE : data <= 8'b00000000 ;
			15'h000024CF : data <= 8'b00000000 ;
			15'h000024D0 : data <= 8'b00000000 ;
			15'h000024D1 : data <= 8'b00000000 ;
			15'h000024D2 : data <= 8'b00000000 ;
			15'h000024D3 : data <= 8'b00000000 ;
			15'h000024D4 : data <= 8'b00000000 ;
			15'h000024D5 : data <= 8'b00000000 ;
			15'h000024D6 : data <= 8'b00000000 ;
			15'h000024D7 : data <= 8'b00000000 ;
			15'h000024D8 : data <= 8'b00000000 ;
			15'h000024D9 : data <= 8'b00000000 ;
			15'h000024DA : data <= 8'b00000000 ;
			15'h000024DB : data <= 8'b00000000 ;
			15'h000024DC : data <= 8'b00000000 ;
			15'h000024DD : data <= 8'b00000000 ;
			15'h000024DE : data <= 8'b00000000 ;
			15'h000024DF : data <= 8'b00000000 ;
			15'h000024E0 : data <= 8'b00000000 ;
			15'h000024E1 : data <= 8'b00000000 ;
			15'h000024E2 : data <= 8'b00000000 ;
			15'h000024E3 : data <= 8'b00000000 ;
			15'h000024E4 : data <= 8'b00000000 ;
			15'h000024E5 : data <= 8'b00000000 ;
			15'h000024E6 : data <= 8'b00000000 ;
			15'h000024E7 : data <= 8'b00000000 ;
			15'h000024E8 : data <= 8'b00000000 ;
			15'h000024E9 : data <= 8'b00000000 ;
			15'h000024EA : data <= 8'b00000000 ;
			15'h000024EB : data <= 8'b00000000 ;
			15'h000024EC : data <= 8'b00000000 ;
			15'h000024ED : data <= 8'b00000000 ;
			15'h000024EE : data <= 8'b00000000 ;
			15'h000024EF : data <= 8'b00000000 ;
			15'h000024F0 : data <= 8'b00000000 ;
			15'h000024F1 : data <= 8'b00000000 ;
			15'h000024F2 : data <= 8'b00000000 ;
			15'h000024F3 : data <= 8'b00000000 ;
			15'h000024F4 : data <= 8'b00000000 ;
			15'h000024F5 : data <= 8'b00000000 ;
			15'h000024F6 : data <= 8'b00000000 ;
			15'h000024F7 : data <= 8'b00000000 ;
			15'h000024F8 : data <= 8'b00000000 ;
			15'h000024F9 : data <= 8'b00000000 ;
			15'h000024FA : data <= 8'b00000000 ;
			15'h000024FB : data <= 8'b00000000 ;
			15'h000024FC : data <= 8'b00000000 ;
			15'h000024FD : data <= 8'b00000000 ;
			15'h000024FE : data <= 8'b00000000 ;
			15'h000024FF : data <= 8'b00000000 ;
			15'h00002500 : data <= 8'b00000000 ;
			15'h00002501 : data <= 8'b00000000 ;
			15'h00002502 : data <= 8'b00000000 ;
			15'h00002503 : data <= 8'b00000000 ;
			15'h00002504 : data <= 8'b00000000 ;
			15'h00002505 : data <= 8'b00000000 ;
			15'h00002506 : data <= 8'b00000000 ;
			15'h00002507 : data <= 8'b00000000 ;
			15'h00002508 : data <= 8'b00000000 ;
			15'h00002509 : data <= 8'b00000000 ;
			15'h0000250A : data <= 8'b00000000 ;
			15'h0000250B : data <= 8'b00000000 ;
			15'h0000250C : data <= 8'b00000000 ;
			15'h0000250D : data <= 8'b00000000 ;
			15'h0000250E : data <= 8'b00000000 ;
			15'h0000250F : data <= 8'b00000000 ;
			15'h00002510 : data <= 8'b00000000 ;
			15'h00002511 : data <= 8'b00000000 ;
			15'h00002512 : data <= 8'b00000000 ;
			15'h00002513 : data <= 8'b00000000 ;
			15'h00002514 : data <= 8'b00000000 ;
			15'h00002515 : data <= 8'b00000000 ;
			15'h00002516 : data <= 8'b00000000 ;
			15'h00002517 : data <= 8'b00000000 ;
			15'h00002518 : data <= 8'b00000000 ;
			15'h00002519 : data <= 8'b00000000 ;
			15'h0000251A : data <= 8'b00000000 ;
			15'h0000251B : data <= 8'b00000000 ;
			15'h0000251C : data <= 8'b00000000 ;
			15'h0000251D : data <= 8'b00000000 ;
			15'h0000251E : data <= 8'b00000000 ;
			15'h0000251F : data <= 8'b00000000 ;
			15'h00002520 : data <= 8'b00000000 ;
			15'h00002521 : data <= 8'b00000000 ;
			15'h00002522 : data <= 8'b00000000 ;
			15'h00002523 : data <= 8'b00000000 ;
			15'h00002524 : data <= 8'b00000000 ;
			15'h00002525 : data <= 8'b00000000 ;
			15'h00002526 : data <= 8'b00000000 ;
			15'h00002527 : data <= 8'b00000000 ;
			15'h00002528 : data <= 8'b00000000 ;
			15'h00002529 : data <= 8'b00000000 ;
			15'h0000252A : data <= 8'b00000000 ;
			15'h0000252B : data <= 8'b00000000 ;
			15'h0000252C : data <= 8'b00000000 ;
			15'h0000252D : data <= 8'b00000000 ;
			15'h0000252E : data <= 8'b00000000 ;
			15'h0000252F : data <= 8'b00000000 ;
			15'h00002530 : data <= 8'b00000000 ;
			15'h00002531 : data <= 8'b00000000 ;
			15'h00002532 : data <= 8'b00000000 ;
			15'h00002533 : data <= 8'b00000000 ;
			15'h00002534 : data <= 8'b00000000 ;
			15'h00002535 : data <= 8'b00000000 ;
			15'h00002536 : data <= 8'b00000000 ;
			15'h00002537 : data <= 8'b00000000 ;
			15'h00002538 : data <= 8'b00000000 ;
			15'h00002539 : data <= 8'b00000000 ;
			15'h0000253A : data <= 8'b00000000 ;
			15'h0000253B : data <= 8'b00000000 ;
			15'h0000253C : data <= 8'b00000000 ;
			15'h0000253D : data <= 8'b00000000 ;
			15'h0000253E : data <= 8'b00000000 ;
			15'h0000253F : data <= 8'b00000000 ;
			15'h00002540 : data <= 8'b00000000 ;
			15'h00002541 : data <= 8'b00000000 ;
			15'h00002542 : data <= 8'b00000000 ;
			15'h00002543 : data <= 8'b00000000 ;
			15'h00002544 : data <= 8'b00000000 ;
			15'h00002545 : data <= 8'b00000000 ;
			15'h00002546 : data <= 8'b00000000 ;
			15'h00002547 : data <= 8'b00000000 ;
			15'h00002548 : data <= 8'b00000000 ;
			15'h00002549 : data <= 8'b00000000 ;
			15'h0000254A : data <= 8'b00000000 ;
			15'h0000254B : data <= 8'b00000000 ;
			15'h0000254C : data <= 8'b00000000 ;
			15'h0000254D : data <= 8'b00000000 ;
			15'h0000254E : data <= 8'b00000000 ;
			15'h0000254F : data <= 8'b00000000 ;
			15'h00002550 : data <= 8'b00000000 ;
			15'h00002551 : data <= 8'b00000000 ;
			15'h00002552 : data <= 8'b00000000 ;
			15'h00002553 : data <= 8'b00000000 ;
			15'h00002554 : data <= 8'b00000000 ;
			15'h00002555 : data <= 8'b00000000 ;
			15'h00002556 : data <= 8'b00000000 ;
			15'h00002557 : data <= 8'b00000000 ;
			15'h00002558 : data <= 8'b00000000 ;
			15'h00002559 : data <= 8'b00000000 ;
			15'h0000255A : data <= 8'b00000000 ;
			15'h0000255B : data <= 8'b00000000 ;
			15'h0000255C : data <= 8'b00000000 ;
			15'h0000255D : data <= 8'b00000000 ;
			15'h0000255E : data <= 8'b00000000 ;
			15'h0000255F : data <= 8'b00000000 ;
			15'h00002560 : data <= 8'b00000000 ;
			15'h00002561 : data <= 8'b00000000 ;
			15'h00002562 : data <= 8'b00000000 ;
			15'h00002563 : data <= 8'b00000000 ;
			15'h00002564 : data <= 8'b00000000 ;
			15'h00002565 : data <= 8'b00000000 ;
			15'h00002566 : data <= 8'b00000000 ;
			15'h00002567 : data <= 8'b00000000 ;
			15'h00002568 : data <= 8'b00000000 ;
			15'h00002569 : data <= 8'b00000000 ;
			15'h0000256A : data <= 8'b00000000 ;
			15'h0000256B : data <= 8'b00000000 ;
			15'h0000256C : data <= 8'b00000000 ;
			15'h0000256D : data <= 8'b00000000 ;
			15'h0000256E : data <= 8'b00000000 ;
			15'h0000256F : data <= 8'b00000000 ;
			15'h00002570 : data <= 8'b00000000 ;
			15'h00002571 : data <= 8'b00000000 ;
			15'h00002572 : data <= 8'b00000000 ;
			15'h00002573 : data <= 8'b00000000 ;
			15'h00002574 : data <= 8'b00000000 ;
			15'h00002575 : data <= 8'b00000000 ;
			15'h00002576 : data <= 8'b00000000 ;
			15'h00002577 : data <= 8'b00000000 ;
			15'h00002578 : data <= 8'b00000000 ;
			15'h00002579 : data <= 8'b00000000 ;
			15'h0000257A : data <= 8'b00000000 ;
			15'h0000257B : data <= 8'b00000000 ;
			15'h0000257C : data <= 8'b00000000 ;
			15'h0000257D : data <= 8'b00000000 ;
			15'h0000257E : data <= 8'b00000000 ;
			15'h0000257F : data <= 8'b00000000 ;
			15'h00002580 : data <= 8'b00000000 ;
			15'h00002581 : data <= 8'b00000000 ;
			15'h00002582 : data <= 8'b00000000 ;
			15'h00002583 : data <= 8'b00000000 ;
			15'h00002584 : data <= 8'b00000000 ;
			15'h00002585 : data <= 8'b00000000 ;
			15'h00002586 : data <= 8'b00000000 ;
			15'h00002587 : data <= 8'b00000000 ;
			15'h00002588 : data <= 8'b00000000 ;
			15'h00002589 : data <= 8'b00000000 ;
			15'h0000258A : data <= 8'b00000000 ;
			15'h0000258B : data <= 8'b00000000 ;
			15'h0000258C : data <= 8'b00000000 ;
			15'h0000258D : data <= 8'b00000000 ;
			15'h0000258E : data <= 8'b00000000 ;
			15'h0000258F : data <= 8'b00000000 ;
			15'h00002590 : data <= 8'b00000000 ;
			15'h00002591 : data <= 8'b00000000 ;
			15'h00002592 : data <= 8'b00000000 ;
			15'h00002593 : data <= 8'b00000000 ;
			15'h00002594 : data <= 8'b00000000 ;
			15'h00002595 : data <= 8'b00000000 ;
			15'h00002596 : data <= 8'b00000000 ;
			15'h00002597 : data <= 8'b00000000 ;
			15'h00002598 : data <= 8'b00000000 ;
			15'h00002599 : data <= 8'b00000000 ;
			15'h0000259A : data <= 8'b00000000 ;
			15'h0000259B : data <= 8'b00000000 ;
			15'h0000259C : data <= 8'b00000000 ;
			15'h0000259D : data <= 8'b00000000 ;
			15'h0000259E : data <= 8'b00000000 ;
			15'h0000259F : data <= 8'b00000000 ;
			15'h000025A0 : data <= 8'b00000000 ;
			15'h000025A1 : data <= 8'b00000000 ;
			15'h000025A2 : data <= 8'b00000000 ;
			15'h000025A3 : data <= 8'b00000000 ;
			15'h000025A4 : data <= 8'b00000000 ;
			15'h000025A5 : data <= 8'b00000000 ;
			15'h000025A6 : data <= 8'b00000000 ;
			15'h000025A7 : data <= 8'b00000000 ;
			15'h000025A8 : data <= 8'b00000000 ;
			15'h000025A9 : data <= 8'b00000000 ;
			15'h000025AA : data <= 8'b00000000 ;
			15'h000025AB : data <= 8'b00000000 ;
			15'h000025AC : data <= 8'b00000000 ;
			15'h000025AD : data <= 8'b00000000 ;
			15'h000025AE : data <= 8'b00000000 ;
			15'h000025AF : data <= 8'b00000000 ;
			15'h000025B0 : data <= 8'b00000000 ;
			15'h000025B1 : data <= 8'b00000000 ;
			15'h000025B2 : data <= 8'b00000000 ;
			15'h000025B3 : data <= 8'b00000000 ;
			15'h000025B4 : data <= 8'b00000000 ;
			15'h000025B5 : data <= 8'b00000000 ;
			15'h000025B6 : data <= 8'b00000000 ;
			15'h000025B7 : data <= 8'b00000000 ;
			15'h000025B8 : data <= 8'b00000000 ;
			15'h000025B9 : data <= 8'b00000000 ;
			15'h000025BA : data <= 8'b00000000 ;
			15'h000025BB : data <= 8'b00000000 ;
			15'h000025BC : data <= 8'b00000000 ;
			15'h000025BD : data <= 8'b00000000 ;
			15'h000025BE : data <= 8'b00000000 ;
			15'h000025BF : data <= 8'b00000000 ;
			15'h000025C0 : data <= 8'b00000000 ;
			15'h000025C1 : data <= 8'b00000000 ;
			15'h000025C2 : data <= 8'b00000000 ;
			15'h000025C3 : data <= 8'b00000000 ;
			15'h000025C4 : data <= 8'b00000000 ;
			15'h000025C5 : data <= 8'b00000000 ;
			15'h000025C6 : data <= 8'b00000000 ;
			15'h000025C7 : data <= 8'b00000000 ;
			15'h000025C8 : data <= 8'b00000000 ;
			15'h000025C9 : data <= 8'b00000000 ;
			15'h000025CA : data <= 8'b00000000 ;
			15'h000025CB : data <= 8'b00000000 ;
			15'h000025CC : data <= 8'b00000000 ;
			15'h000025CD : data <= 8'b00000000 ;
			15'h000025CE : data <= 8'b00000000 ;
			15'h000025CF : data <= 8'b00000000 ;
			15'h000025D0 : data <= 8'b00000000 ;
			15'h000025D1 : data <= 8'b00000000 ;
			15'h000025D2 : data <= 8'b00000000 ;
			15'h000025D3 : data <= 8'b00000000 ;
			15'h000025D4 : data <= 8'b00000000 ;
			15'h000025D5 : data <= 8'b00000000 ;
			15'h000025D6 : data <= 8'b00000000 ;
			15'h000025D7 : data <= 8'b00000000 ;
			15'h000025D8 : data <= 8'b00000000 ;
			15'h000025D9 : data <= 8'b00000000 ;
			15'h000025DA : data <= 8'b00000000 ;
			15'h000025DB : data <= 8'b00000000 ;
			15'h000025DC : data <= 8'b00000000 ;
			15'h000025DD : data <= 8'b00000000 ;
			15'h000025DE : data <= 8'b00000000 ;
			15'h000025DF : data <= 8'b00000000 ;
			15'h000025E0 : data <= 8'b00000000 ;
			15'h000025E1 : data <= 8'b00000000 ;
			15'h000025E2 : data <= 8'b00000000 ;
			15'h000025E3 : data <= 8'b00000000 ;
			15'h000025E4 : data <= 8'b00000000 ;
			15'h000025E5 : data <= 8'b00000000 ;
			15'h000025E6 : data <= 8'b00000000 ;
			15'h000025E7 : data <= 8'b00000000 ;
			15'h000025E8 : data <= 8'b00000000 ;
			15'h000025E9 : data <= 8'b00000000 ;
			15'h000025EA : data <= 8'b00000000 ;
			15'h000025EB : data <= 8'b00000000 ;
			15'h000025EC : data <= 8'b00000000 ;
			15'h000025ED : data <= 8'b00000000 ;
			15'h000025EE : data <= 8'b00000000 ;
			15'h000025EF : data <= 8'b00000000 ;
			15'h000025F0 : data <= 8'b00000000 ;
			15'h000025F1 : data <= 8'b00000000 ;
			15'h000025F2 : data <= 8'b00000000 ;
			15'h000025F3 : data <= 8'b00000000 ;
			15'h000025F4 : data <= 8'b00000000 ;
			15'h000025F5 : data <= 8'b00000000 ;
			15'h000025F6 : data <= 8'b00000000 ;
			15'h000025F7 : data <= 8'b00000000 ;
			15'h000025F8 : data <= 8'b00000000 ;
			15'h000025F9 : data <= 8'b00000000 ;
			15'h000025FA : data <= 8'b00000000 ;
			15'h000025FB : data <= 8'b00000000 ;
			15'h000025FC : data <= 8'b00000000 ;
			15'h000025FD : data <= 8'b00000000 ;
			15'h000025FE : data <= 8'b00000000 ;
			15'h000025FF : data <= 8'b00000000 ;
			15'h00002600 : data <= 8'b00000000 ;
			15'h00002601 : data <= 8'b00000000 ;
			15'h00002602 : data <= 8'b00000000 ;
			15'h00002603 : data <= 8'b00000000 ;
			15'h00002604 : data <= 8'b00000000 ;
			15'h00002605 : data <= 8'b00000000 ;
			15'h00002606 : data <= 8'b00000000 ;
			15'h00002607 : data <= 8'b00000000 ;
			15'h00002608 : data <= 8'b00000000 ;
			15'h00002609 : data <= 8'b00000000 ;
			15'h0000260A : data <= 8'b00000000 ;
			15'h0000260B : data <= 8'b00000000 ;
			15'h0000260C : data <= 8'b00000000 ;
			15'h0000260D : data <= 8'b00000000 ;
			15'h0000260E : data <= 8'b00000000 ;
			15'h0000260F : data <= 8'b00000000 ;
			15'h00002610 : data <= 8'b00000000 ;
			15'h00002611 : data <= 8'b00000000 ;
			15'h00002612 : data <= 8'b00000000 ;
			15'h00002613 : data <= 8'b00000000 ;
			15'h00002614 : data <= 8'b00000000 ;
			15'h00002615 : data <= 8'b00000000 ;
			15'h00002616 : data <= 8'b00000000 ;
			15'h00002617 : data <= 8'b00000000 ;
			15'h00002618 : data <= 8'b00000000 ;
			15'h00002619 : data <= 8'b00000000 ;
			15'h0000261A : data <= 8'b00000000 ;
			15'h0000261B : data <= 8'b00000000 ;
			15'h0000261C : data <= 8'b00000000 ;
			15'h0000261D : data <= 8'b00000000 ;
			15'h0000261E : data <= 8'b00000000 ;
			15'h0000261F : data <= 8'b00000000 ;
			15'h00002620 : data <= 8'b00000000 ;
			15'h00002621 : data <= 8'b00000000 ;
			15'h00002622 : data <= 8'b00000000 ;
			15'h00002623 : data <= 8'b00000000 ;
			15'h00002624 : data <= 8'b00000000 ;
			15'h00002625 : data <= 8'b00000000 ;
			15'h00002626 : data <= 8'b00000000 ;
			15'h00002627 : data <= 8'b00000000 ;
			15'h00002628 : data <= 8'b00000000 ;
			15'h00002629 : data <= 8'b00000000 ;
			15'h0000262A : data <= 8'b00000000 ;
			15'h0000262B : data <= 8'b00000000 ;
			15'h0000262C : data <= 8'b00000000 ;
			15'h0000262D : data <= 8'b00000000 ;
			15'h0000262E : data <= 8'b00000000 ;
			15'h0000262F : data <= 8'b00000000 ;
			15'h00002630 : data <= 8'b00000000 ;
			15'h00002631 : data <= 8'b00000000 ;
			15'h00002632 : data <= 8'b00000000 ;
			15'h00002633 : data <= 8'b00000000 ;
			15'h00002634 : data <= 8'b00000000 ;
			15'h00002635 : data <= 8'b00000000 ;
			15'h00002636 : data <= 8'b00000000 ;
			15'h00002637 : data <= 8'b00000000 ;
			15'h00002638 : data <= 8'b00000000 ;
			15'h00002639 : data <= 8'b00000000 ;
			15'h0000263A : data <= 8'b00000000 ;
			15'h0000263B : data <= 8'b00000000 ;
			15'h0000263C : data <= 8'b00000000 ;
			15'h0000263D : data <= 8'b00000000 ;
			15'h0000263E : data <= 8'b00000000 ;
			15'h0000263F : data <= 8'b00000000 ;
			15'h00002640 : data <= 8'b00000000 ;
			15'h00002641 : data <= 8'b00000000 ;
			15'h00002642 : data <= 8'b00000000 ;
			15'h00002643 : data <= 8'b00000000 ;
			15'h00002644 : data <= 8'b00000000 ;
			15'h00002645 : data <= 8'b00000000 ;
			15'h00002646 : data <= 8'b00000000 ;
			15'h00002647 : data <= 8'b00000000 ;
			15'h00002648 : data <= 8'b00000000 ;
			15'h00002649 : data <= 8'b00000000 ;
			15'h0000264A : data <= 8'b00000000 ;
			15'h0000264B : data <= 8'b00000000 ;
			15'h0000264C : data <= 8'b00000000 ;
			15'h0000264D : data <= 8'b00000000 ;
			15'h0000264E : data <= 8'b00000000 ;
			15'h0000264F : data <= 8'b00000000 ;
			15'h00002650 : data <= 8'b00000000 ;
			15'h00002651 : data <= 8'b00000000 ;
			15'h00002652 : data <= 8'b00000000 ;
			15'h00002653 : data <= 8'b00000000 ;
			15'h00002654 : data <= 8'b00000000 ;
			15'h00002655 : data <= 8'b00000000 ;
			15'h00002656 : data <= 8'b00000000 ;
			15'h00002657 : data <= 8'b00000000 ;
			15'h00002658 : data <= 8'b00000000 ;
			15'h00002659 : data <= 8'b00000000 ;
			15'h0000265A : data <= 8'b00000000 ;
			15'h0000265B : data <= 8'b00000000 ;
			15'h0000265C : data <= 8'b00000000 ;
			15'h0000265D : data <= 8'b00000000 ;
			15'h0000265E : data <= 8'b00000000 ;
			15'h0000265F : data <= 8'b00000000 ;
			15'h00002660 : data <= 8'b00000000 ;
			15'h00002661 : data <= 8'b00000000 ;
			15'h00002662 : data <= 8'b00000000 ;
			15'h00002663 : data <= 8'b00000000 ;
			15'h00002664 : data <= 8'b00000000 ;
			15'h00002665 : data <= 8'b00000000 ;
			15'h00002666 : data <= 8'b00000000 ;
			15'h00002667 : data <= 8'b00000000 ;
			15'h00002668 : data <= 8'b00000000 ;
			15'h00002669 : data <= 8'b00000000 ;
			15'h0000266A : data <= 8'b00000000 ;
			15'h0000266B : data <= 8'b00000000 ;
			15'h0000266C : data <= 8'b00000000 ;
			15'h0000266D : data <= 8'b00000000 ;
			15'h0000266E : data <= 8'b00000000 ;
			15'h0000266F : data <= 8'b00000000 ;
			15'h00002670 : data <= 8'b00000000 ;
			15'h00002671 : data <= 8'b00000000 ;
			15'h00002672 : data <= 8'b00000000 ;
			15'h00002673 : data <= 8'b00000000 ;
			15'h00002674 : data <= 8'b00000000 ;
			15'h00002675 : data <= 8'b00000000 ;
			15'h00002676 : data <= 8'b00000000 ;
			15'h00002677 : data <= 8'b00000000 ;
			15'h00002678 : data <= 8'b00000000 ;
			15'h00002679 : data <= 8'b00000000 ;
			15'h0000267A : data <= 8'b00000000 ;
			15'h0000267B : data <= 8'b00000000 ;
			15'h0000267C : data <= 8'b00000000 ;
			15'h0000267D : data <= 8'b00000000 ;
			15'h0000267E : data <= 8'b00000000 ;
			15'h0000267F : data <= 8'b00000000 ;
			15'h00002680 : data <= 8'b00000000 ;
			15'h00002681 : data <= 8'b00000000 ;
			15'h00002682 : data <= 8'b00000000 ;
			15'h00002683 : data <= 8'b00000000 ;
			15'h00002684 : data <= 8'b00000000 ;
			15'h00002685 : data <= 8'b00000000 ;
			15'h00002686 : data <= 8'b00000000 ;
			15'h00002687 : data <= 8'b00000000 ;
			15'h00002688 : data <= 8'b00000000 ;
			15'h00002689 : data <= 8'b00000000 ;
			15'h0000268A : data <= 8'b00000000 ;
			15'h0000268B : data <= 8'b00000000 ;
			15'h0000268C : data <= 8'b00000000 ;
			15'h0000268D : data <= 8'b00000000 ;
			15'h0000268E : data <= 8'b00000000 ;
			15'h0000268F : data <= 8'b00000000 ;
			15'h00002690 : data <= 8'b00000000 ;
			15'h00002691 : data <= 8'b00000000 ;
			15'h00002692 : data <= 8'b00000000 ;
			15'h00002693 : data <= 8'b00000000 ;
			15'h00002694 : data <= 8'b00000000 ;
			15'h00002695 : data <= 8'b00000000 ;
			15'h00002696 : data <= 8'b00000000 ;
			15'h00002697 : data <= 8'b00000000 ;
			15'h00002698 : data <= 8'b00000000 ;
			15'h00002699 : data <= 8'b00000000 ;
			15'h0000269A : data <= 8'b00000000 ;
			15'h0000269B : data <= 8'b00000000 ;
			15'h0000269C : data <= 8'b00000000 ;
			15'h0000269D : data <= 8'b00000000 ;
			15'h0000269E : data <= 8'b00000000 ;
			15'h0000269F : data <= 8'b00000000 ;
			15'h000026A0 : data <= 8'b00000000 ;
			15'h000026A1 : data <= 8'b00000000 ;
			15'h000026A2 : data <= 8'b00000000 ;
			15'h000026A3 : data <= 8'b00000000 ;
			15'h000026A4 : data <= 8'b00000000 ;
			15'h000026A5 : data <= 8'b00000000 ;
			15'h000026A6 : data <= 8'b00000000 ;
			15'h000026A7 : data <= 8'b00000000 ;
			15'h000026A8 : data <= 8'b00000000 ;
			15'h000026A9 : data <= 8'b00000000 ;
			15'h000026AA : data <= 8'b00000000 ;
			15'h000026AB : data <= 8'b00000000 ;
			15'h000026AC : data <= 8'b00000000 ;
			15'h000026AD : data <= 8'b00000000 ;
			15'h000026AE : data <= 8'b00000000 ;
			15'h000026AF : data <= 8'b00000000 ;
			15'h000026B0 : data <= 8'b00000000 ;
			15'h000026B1 : data <= 8'b00000000 ;
			15'h000026B2 : data <= 8'b00000000 ;
			15'h000026B3 : data <= 8'b00000000 ;
			15'h000026B4 : data <= 8'b00000000 ;
			15'h000026B5 : data <= 8'b00000000 ;
			15'h000026B6 : data <= 8'b00000000 ;
			15'h000026B7 : data <= 8'b00000000 ;
			15'h000026B8 : data <= 8'b00000000 ;
			15'h000026B9 : data <= 8'b00000000 ;
			15'h000026BA : data <= 8'b00000000 ;
			15'h000026BB : data <= 8'b00000000 ;
			15'h000026BC : data <= 8'b00000000 ;
			15'h000026BD : data <= 8'b00000000 ;
			15'h000026BE : data <= 8'b00000000 ;
			15'h000026BF : data <= 8'b00000000 ;
			15'h000026C0 : data <= 8'b00000000 ;
			15'h000026C1 : data <= 8'b00000000 ;
			15'h000026C2 : data <= 8'b00000000 ;
			15'h000026C3 : data <= 8'b00000000 ;
			15'h000026C4 : data <= 8'b00000000 ;
			15'h000026C5 : data <= 8'b00000000 ;
			15'h000026C6 : data <= 8'b00000000 ;
			15'h000026C7 : data <= 8'b00000000 ;
			15'h000026C8 : data <= 8'b00000000 ;
			15'h000026C9 : data <= 8'b00000000 ;
			15'h000026CA : data <= 8'b00000000 ;
			15'h000026CB : data <= 8'b00000000 ;
			15'h000026CC : data <= 8'b00000000 ;
			15'h000026CD : data <= 8'b00000000 ;
			15'h000026CE : data <= 8'b00000000 ;
			15'h000026CF : data <= 8'b00000000 ;
			15'h000026D0 : data <= 8'b00000000 ;
			15'h000026D1 : data <= 8'b00000000 ;
			15'h000026D2 : data <= 8'b00000000 ;
			15'h000026D3 : data <= 8'b00000000 ;
			15'h000026D4 : data <= 8'b00000000 ;
			15'h000026D5 : data <= 8'b00000000 ;
			15'h000026D6 : data <= 8'b00000000 ;
			15'h000026D7 : data <= 8'b00000000 ;
			15'h000026D8 : data <= 8'b00000000 ;
			15'h000026D9 : data <= 8'b00000000 ;
			15'h000026DA : data <= 8'b00000000 ;
			15'h000026DB : data <= 8'b00000000 ;
			15'h000026DC : data <= 8'b00000000 ;
			15'h000026DD : data <= 8'b00000000 ;
			15'h000026DE : data <= 8'b00000000 ;
			15'h000026DF : data <= 8'b00000000 ;
			15'h000026E0 : data <= 8'b00000000 ;
			15'h000026E1 : data <= 8'b00000000 ;
			15'h000026E2 : data <= 8'b00000000 ;
			15'h000026E3 : data <= 8'b00000000 ;
			15'h000026E4 : data <= 8'b00000000 ;
			15'h000026E5 : data <= 8'b00000000 ;
			15'h000026E6 : data <= 8'b00000000 ;
			15'h000026E7 : data <= 8'b00000000 ;
			15'h000026E8 : data <= 8'b00000000 ;
			15'h000026E9 : data <= 8'b00000000 ;
			15'h000026EA : data <= 8'b00000000 ;
			15'h000026EB : data <= 8'b00000000 ;
			15'h000026EC : data <= 8'b00000000 ;
			15'h000026ED : data <= 8'b00000000 ;
			15'h000026EE : data <= 8'b00000000 ;
			15'h000026EF : data <= 8'b00000000 ;
			15'h000026F0 : data <= 8'b00000000 ;
			15'h000026F1 : data <= 8'b00000000 ;
			15'h000026F2 : data <= 8'b00000000 ;
			15'h000026F3 : data <= 8'b00000000 ;
			15'h000026F4 : data <= 8'b00000000 ;
			15'h000026F5 : data <= 8'b00000000 ;
			15'h000026F6 : data <= 8'b00000000 ;
			15'h000026F7 : data <= 8'b00000000 ;
			15'h000026F8 : data <= 8'b00000000 ;
			15'h000026F9 : data <= 8'b00000000 ;
			15'h000026FA : data <= 8'b00000000 ;
			15'h000026FB : data <= 8'b00000000 ;
			15'h000026FC : data <= 8'b00000000 ;
			15'h000026FD : data <= 8'b00000000 ;
			15'h000026FE : data <= 8'b00000000 ;
			15'h000026FF : data <= 8'b00000000 ;
			15'h00002700 : data <= 8'b00000000 ;
			15'h00002701 : data <= 8'b00000000 ;
			15'h00002702 : data <= 8'b00000000 ;
			15'h00002703 : data <= 8'b00000000 ;
			15'h00002704 : data <= 8'b00000000 ;
			15'h00002705 : data <= 8'b00000000 ;
			15'h00002706 : data <= 8'b00000000 ;
			15'h00002707 : data <= 8'b00000000 ;
			15'h00002708 : data <= 8'b00000000 ;
			15'h00002709 : data <= 8'b00000000 ;
			15'h0000270A : data <= 8'b00000000 ;
			15'h0000270B : data <= 8'b00000000 ;
			15'h0000270C : data <= 8'b00000000 ;
			15'h0000270D : data <= 8'b00000000 ;
			15'h0000270E : data <= 8'b00000000 ;
			15'h0000270F : data <= 8'b00000000 ;
			15'h00002710 : data <= 8'b00000000 ;
			15'h00002711 : data <= 8'b00000000 ;
			15'h00002712 : data <= 8'b00000000 ;
			15'h00002713 : data <= 8'b00000000 ;
			15'h00002714 : data <= 8'b00000000 ;
			15'h00002715 : data <= 8'b00000000 ;
			15'h00002716 : data <= 8'b00000000 ;
			15'h00002717 : data <= 8'b00000000 ;
			15'h00002718 : data <= 8'b00000000 ;
			15'h00002719 : data <= 8'b00000000 ;
			15'h0000271A : data <= 8'b00000000 ;
			15'h0000271B : data <= 8'b00000000 ;
			15'h0000271C : data <= 8'b00000000 ;
			15'h0000271D : data <= 8'b00000000 ;
			15'h0000271E : data <= 8'b00000000 ;
			15'h0000271F : data <= 8'b00000000 ;
			15'h00002720 : data <= 8'b00000000 ;
			15'h00002721 : data <= 8'b00000000 ;
			15'h00002722 : data <= 8'b00000000 ;
			15'h00002723 : data <= 8'b00000000 ;
			15'h00002724 : data <= 8'b00000000 ;
			15'h00002725 : data <= 8'b00000000 ;
			15'h00002726 : data <= 8'b00000000 ;
			15'h00002727 : data <= 8'b00000000 ;
			15'h00002728 : data <= 8'b00000000 ;
			15'h00002729 : data <= 8'b00000000 ;
			15'h0000272A : data <= 8'b00000000 ;
			15'h0000272B : data <= 8'b00000000 ;
			15'h0000272C : data <= 8'b00000000 ;
			15'h0000272D : data <= 8'b00000000 ;
			15'h0000272E : data <= 8'b00000000 ;
			15'h0000272F : data <= 8'b00000000 ;
			15'h00002730 : data <= 8'b00000000 ;
			15'h00002731 : data <= 8'b00000000 ;
			15'h00002732 : data <= 8'b00000000 ;
			15'h00002733 : data <= 8'b00000000 ;
			15'h00002734 : data <= 8'b00000000 ;
			15'h00002735 : data <= 8'b00000000 ;
			15'h00002736 : data <= 8'b00000000 ;
			15'h00002737 : data <= 8'b00000000 ;
			15'h00002738 : data <= 8'b00000000 ;
			15'h00002739 : data <= 8'b00000000 ;
			15'h0000273A : data <= 8'b00000000 ;
			15'h0000273B : data <= 8'b00000000 ;
			15'h0000273C : data <= 8'b00000000 ;
			15'h0000273D : data <= 8'b00000000 ;
			15'h0000273E : data <= 8'b00000000 ;
			15'h0000273F : data <= 8'b00000000 ;
			15'h00002740 : data <= 8'b00000000 ;
			15'h00002741 : data <= 8'b00000000 ;
			15'h00002742 : data <= 8'b00000000 ;
			15'h00002743 : data <= 8'b00000000 ;
			15'h00002744 : data <= 8'b00000000 ;
			15'h00002745 : data <= 8'b00000000 ;
			15'h00002746 : data <= 8'b00000000 ;
			15'h00002747 : data <= 8'b00000000 ;
			15'h00002748 : data <= 8'b00000000 ;
			15'h00002749 : data <= 8'b00000000 ;
			15'h0000274A : data <= 8'b00000000 ;
			15'h0000274B : data <= 8'b00000000 ;
			15'h0000274C : data <= 8'b00000000 ;
			15'h0000274D : data <= 8'b00000000 ;
			15'h0000274E : data <= 8'b00000000 ;
			15'h0000274F : data <= 8'b00000000 ;
			15'h00002750 : data <= 8'b00000000 ;
			15'h00002751 : data <= 8'b00000000 ;
			15'h00002752 : data <= 8'b00000000 ;
			15'h00002753 : data <= 8'b00000000 ;
			15'h00002754 : data <= 8'b00000000 ;
			15'h00002755 : data <= 8'b00000000 ;
			15'h00002756 : data <= 8'b00000000 ;
			15'h00002757 : data <= 8'b00000000 ;
			15'h00002758 : data <= 8'b00000000 ;
			15'h00002759 : data <= 8'b00000000 ;
			15'h0000275A : data <= 8'b00000000 ;
			15'h0000275B : data <= 8'b00000000 ;
			15'h0000275C : data <= 8'b00000000 ;
			15'h0000275D : data <= 8'b00000000 ;
			15'h0000275E : data <= 8'b00000000 ;
			15'h0000275F : data <= 8'b00000000 ;
			15'h00002760 : data <= 8'b00000000 ;
			15'h00002761 : data <= 8'b00000000 ;
			15'h00002762 : data <= 8'b00000000 ;
			15'h00002763 : data <= 8'b00000000 ;
			15'h00002764 : data <= 8'b00000000 ;
			15'h00002765 : data <= 8'b00000000 ;
			15'h00002766 : data <= 8'b00000000 ;
			15'h00002767 : data <= 8'b00000000 ;
			15'h00002768 : data <= 8'b00000000 ;
			15'h00002769 : data <= 8'b00000000 ;
			15'h0000276A : data <= 8'b00000000 ;
			15'h0000276B : data <= 8'b00000000 ;
			15'h0000276C : data <= 8'b00000000 ;
			15'h0000276D : data <= 8'b00000000 ;
			15'h0000276E : data <= 8'b00000000 ;
			15'h0000276F : data <= 8'b00000000 ;
			15'h00002770 : data <= 8'b00000000 ;
			15'h00002771 : data <= 8'b00000000 ;
			15'h00002772 : data <= 8'b00000000 ;
			15'h00002773 : data <= 8'b00000000 ;
			15'h00002774 : data <= 8'b00000000 ;
			15'h00002775 : data <= 8'b00000000 ;
			15'h00002776 : data <= 8'b00000000 ;
			15'h00002777 : data <= 8'b00000000 ;
			15'h00002778 : data <= 8'b00000000 ;
			15'h00002779 : data <= 8'b00000000 ;
			15'h0000277A : data <= 8'b00000000 ;
			15'h0000277B : data <= 8'b00000000 ;
			15'h0000277C : data <= 8'b00000000 ;
			15'h0000277D : data <= 8'b00000000 ;
			15'h0000277E : data <= 8'b00000000 ;
			15'h0000277F : data <= 8'b00000000 ;
			15'h00002780 : data <= 8'b00000000 ;
			15'h00002781 : data <= 8'b00000000 ;
			15'h00002782 : data <= 8'b00000000 ;
			15'h00002783 : data <= 8'b00000000 ;
			15'h00002784 : data <= 8'b00000000 ;
			15'h00002785 : data <= 8'b00000000 ;
			15'h00002786 : data <= 8'b00000000 ;
			15'h00002787 : data <= 8'b00000000 ;
			15'h00002788 : data <= 8'b00000000 ;
			15'h00002789 : data <= 8'b00000000 ;
			15'h0000278A : data <= 8'b00000000 ;
			15'h0000278B : data <= 8'b00000000 ;
			15'h0000278C : data <= 8'b00000000 ;
			15'h0000278D : data <= 8'b00000000 ;
			15'h0000278E : data <= 8'b00000000 ;
			15'h0000278F : data <= 8'b00000000 ;
			15'h00002790 : data <= 8'b00000000 ;
			15'h00002791 : data <= 8'b00000000 ;
			15'h00002792 : data <= 8'b00000000 ;
			15'h00002793 : data <= 8'b00000000 ;
			15'h00002794 : data <= 8'b00000000 ;
			15'h00002795 : data <= 8'b00000000 ;
			15'h00002796 : data <= 8'b00000000 ;
			15'h00002797 : data <= 8'b00000000 ;
			15'h00002798 : data <= 8'b00000000 ;
			15'h00002799 : data <= 8'b00000000 ;
			15'h0000279A : data <= 8'b00000000 ;
			15'h0000279B : data <= 8'b00000000 ;
			15'h0000279C : data <= 8'b00000000 ;
			15'h0000279D : data <= 8'b00000000 ;
			15'h0000279E : data <= 8'b00000000 ;
			15'h0000279F : data <= 8'b00000000 ;
			15'h000027A0 : data <= 8'b00000000 ;
			15'h000027A1 : data <= 8'b00000000 ;
			15'h000027A2 : data <= 8'b00000000 ;
			15'h000027A3 : data <= 8'b00000000 ;
			15'h000027A4 : data <= 8'b00000000 ;
			15'h000027A5 : data <= 8'b00000000 ;
			15'h000027A6 : data <= 8'b00000000 ;
			15'h000027A7 : data <= 8'b00000000 ;
			15'h000027A8 : data <= 8'b00000000 ;
			15'h000027A9 : data <= 8'b00000000 ;
			15'h000027AA : data <= 8'b00000000 ;
			15'h000027AB : data <= 8'b00000000 ;
			15'h000027AC : data <= 8'b00000000 ;
			15'h000027AD : data <= 8'b00000000 ;
			15'h000027AE : data <= 8'b00000000 ;
			15'h000027AF : data <= 8'b00000000 ;
			15'h000027B0 : data <= 8'b00000000 ;
			15'h000027B1 : data <= 8'b00000000 ;
			15'h000027B2 : data <= 8'b00000000 ;
			15'h000027B3 : data <= 8'b00000000 ;
			15'h000027B4 : data <= 8'b00000000 ;
			15'h000027B5 : data <= 8'b00000000 ;
			15'h000027B6 : data <= 8'b00000000 ;
			15'h000027B7 : data <= 8'b00000000 ;
			15'h000027B8 : data <= 8'b00000000 ;
			15'h000027B9 : data <= 8'b00000000 ;
			15'h000027BA : data <= 8'b00000000 ;
			15'h000027BB : data <= 8'b00000000 ;
			15'h000027BC : data <= 8'b00000000 ;
			15'h000027BD : data <= 8'b00000000 ;
			15'h000027BE : data <= 8'b00000000 ;
			15'h000027BF : data <= 8'b00000000 ;
			15'h000027C0 : data <= 8'b00000000 ;
			15'h000027C1 : data <= 8'b00000000 ;
			15'h000027C2 : data <= 8'b00000000 ;
			15'h000027C3 : data <= 8'b00000000 ;
			15'h000027C4 : data <= 8'b00000000 ;
			15'h000027C5 : data <= 8'b00000000 ;
			15'h000027C6 : data <= 8'b00000000 ;
			15'h000027C7 : data <= 8'b00000000 ;
			15'h000027C8 : data <= 8'b00000000 ;
			15'h000027C9 : data <= 8'b00000000 ;
			15'h000027CA : data <= 8'b00000000 ;
			15'h000027CB : data <= 8'b00000000 ;
			15'h000027CC : data <= 8'b00000000 ;
			15'h000027CD : data <= 8'b00000000 ;
			15'h000027CE : data <= 8'b00000000 ;
			15'h000027CF : data <= 8'b00000000 ;
			15'h000027D0 : data <= 8'b00000000 ;
			15'h000027D1 : data <= 8'b00000000 ;
			15'h000027D2 : data <= 8'b00000000 ;
			15'h000027D3 : data <= 8'b00000000 ;
			15'h000027D4 : data <= 8'b00000000 ;
			15'h000027D5 : data <= 8'b00000000 ;
			15'h000027D6 : data <= 8'b00000000 ;
			15'h000027D7 : data <= 8'b00000000 ;
			15'h000027D8 : data <= 8'b00000000 ;
			15'h000027D9 : data <= 8'b00000000 ;
			15'h000027DA : data <= 8'b00000000 ;
			15'h000027DB : data <= 8'b00000000 ;
			15'h000027DC : data <= 8'b00000000 ;
			15'h000027DD : data <= 8'b00000000 ;
			15'h000027DE : data <= 8'b00000000 ;
			15'h000027DF : data <= 8'b00000000 ;
			15'h000027E0 : data <= 8'b00000000 ;
			15'h000027E1 : data <= 8'b00000000 ;
			15'h000027E2 : data <= 8'b00000000 ;
			15'h000027E3 : data <= 8'b00000000 ;
			15'h000027E4 : data <= 8'b00000000 ;
			15'h000027E5 : data <= 8'b00000000 ;
			15'h000027E6 : data <= 8'b00000000 ;
			15'h000027E7 : data <= 8'b00000000 ;
			15'h000027E8 : data <= 8'b00000000 ;
			15'h000027E9 : data <= 8'b00000000 ;
			15'h000027EA : data <= 8'b00000000 ;
			15'h000027EB : data <= 8'b00000000 ;
			15'h000027EC : data <= 8'b00000000 ;
			15'h000027ED : data <= 8'b00000000 ;
			15'h000027EE : data <= 8'b00000000 ;
			15'h000027EF : data <= 8'b00000000 ;
			15'h000027F0 : data <= 8'b00000000 ;
			15'h000027F1 : data <= 8'b00000000 ;
			15'h000027F2 : data <= 8'b00000000 ;
			15'h000027F3 : data <= 8'b00000000 ;
			15'h000027F4 : data <= 8'b00000000 ;
			15'h000027F5 : data <= 8'b00000000 ;
			15'h000027F6 : data <= 8'b00000000 ;
			15'h000027F7 : data <= 8'b00000000 ;
			15'h000027F8 : data <= 8'b00000000 ;
			15'h000027F9 : data <= 8'b00000000 ;
			15'h000027FA : data <= 8'b00000000 ;
			15'h000027FB : data <= 8'b00000000 ;
			15'h000027FC : data <= 8'b00000000 ;
			15'h000027FD : data <= 8'b00000000 ;
			15'h000027FE : data <= 8'b00000000 ;
			15'h000027FF : data <= 8'b00000000 ;
			15'h00002800 : data <= 8'b00000000 ;
			15'h00002801 : data <= 8'b00000000 ;
			15'h00002802 : data <= 8'b00000000 ;
			15'h00002803 : data <= 8'b00000000 ;
			15'h00002804 : data <= 8'b00000000 ;
			15'h00002805 : data <= 8'b00000000 ;
			15'h00002806 : data <= 8'b00000000 ;
			15'h00002807 : data <= 8'b00000000 ;
			15'h00002808 : data <= 8'b00000000 ;
			15'h00002809 : data <= 8'b00000000 ;
			15'h0000280A : data <= 8'b00000000 ;
			15'h0000280B : data <= 8'b00000000 ;
			15'h0000280C : data <= 8'b00000000 ;
			15'h0000280D : data <= 8'b00000000 ;
			15'h0000280E : data <= 8'b00000000 ;
			15'h0000280F : data <= 8'b00000000 ;
			15'h00002810 : data <= 8'b00000000 ;
			15'h00002811 : data <= 8'b00000000 ;
			15'h00002812 : data <= 8'b00000000 ;
			15'h00002813 : data <= 8'b00000000 ;
			15'h00002814 : data <= 8'b00000000 ;
			15'h00002815 : data <= 8'b00000000 ;
			15'h00002816 : data <= 8'b00000000 ;
			15'h00002817 : data <= 8'b00000000 ;
			15'h00002818 : data <= 8'b00000000 ;
			15'h00002819 : data <= 8'b00000000 ;
			15'h0000281A : data <= 8'b00000000 ;
			15'h0000281B : data <= 8'b00000000 ;
			15'h0000281C : data <= 8'b00000000 ;
			15'h0000281D : data <= 8'b00000000 ;
			15'h0000281E : data <= 8'b00000000 ;
			15'h0000281F : data <= 8'b00000000 ;
			15'h00002820 : data <= 8'b00000000 ;
			15'h00002821 : data <= 8'b00000000 ;
			15'h00002822 : data <= 8'b00000000 ;
			15'h00002823 : data <= 8'b00000000 ;
			15'h00002824 : data <= 8'b00000000 ;
			15'h00002825 : data <= 8'b00000000 ;
			15'h00002826 : data <= 8'b00000000 ;
			15'h00002827 : data <= 8'b00000000 ;
			15'h00002828 : data <= 8'b00000000 ;
			15'h00002829 : data <= 8'b00000000 ;
			15'h0000282A : data <= 8'b00000000 ;
			15'h0000282B : data <= 8'b00000000 ;
			15'h0000282C : data <= 8'b00000000 ;
			15'h0000282D : data <= 8'b00000000 ;
			15'h0000282E : data <= 8'b00000000 ;
			15'h0000282F : data <= 8'b00000000 ;
			15'h00002830 : data <= 8'b00000000 ;
			15'h00002831 : data <= 8'b00000000 ;
			15'h00002832 : data <= 8'b00000000 ;
			15'h00002833 : data <= 8'b00000000 ;
			15'h00002834 : data <= 8'b00000000 ;
			15'h00002835 : data <= 8'b00000000 ;
			15'h00002836 : data <= 8'b00000000 ;
			15'h00002837 : data <= 8'b00000000 ;
			15'h00002838 : data <= 8'b00000000 ;
			15'h00002839 : data <= 8'b00000000 ;
			15'h0000283A : data <= 8'b00000000 ;
			15'h0000283B : data <= 8'b00000000 ;
			15'h0000283C : data <= 8'b00000000 ;
			15'h0000283D : data <= 8'b00000000 ;
			15'h0000283E : data <= 8'b00000000 ;
			15'h0000283F : data <= 8'b00000000 ;
			15'h00002840 : data <= 8'b00000000 ;
			15'h00002841 : data <= 8'b00000000 ;
			15'h00002842 : data <= 8'b00000000 ;
			15'h00002843 : data <= 8'b00000000 ;
			15'h00002844 : data <= 8'b00000000 ;
			15'h00002845 : data <= 8'b00000000 ;
			15'h00002846 : data <= 8'b00000000 ;
			15'h00002847 : data <= 8'b00000000 ;
			15'h00002848 : data <= 8'b00000000 ;
			15'h00002849 : data <= 8'b00000000 ;
			15'h0000284A : data <= 8'b00000000 ;
			15'h0000284B : data <= 8'b00000000 ;
			15'h0000284C : data <= 8'b00000000 ;
			15'h0000284D : data <= 8'b00000000 ;
			15'h0000284E : data <= 8'b00000000 ;
			15'h0000284F : data <= 8'b00000000 ;
			15'h00002850 : data <= 8'b00000000 ;
			15'h00002851 : data <= 8'b00000000 ;
			15'h00002852 : data <= 8'b00000000 ;
			15'h00002853 : data <= 8'b00000000 ;
			15'h00002854 : data <= 8'b00000000 ;
			15'h00002855 : data <= 8'b00000000 ;
			15'h00002856 : data <= 8'b00000000 ;
			15'h00002857 : data <= 8'b00000000 ;
			15'h00002858 : data <= 8'b00000000 ;
			15'h00002859 : data <= 8'b00000000 ;
			15'h0000285A : data <= 8'b00000000 ;
			15'h0000285B : data <= 8'b00000000 ;
			15'h0000285C : data <= 8'b00000000 ;
			15'h0000285D : data <= 8'b00000000 ;
			15'h0000285E : data <= 8'b00000000 ;
			15'h0000285F : data <= 8'b00000000 ;
			15'h00002860 : data <= 8'b00000000 ;
			15'h00002861 : data <= 8'b00000000 ;
			15'h00002862 : data <= 8'b00000000 ;
			15'h00002863 : data <= 8'b00000000 ;
			15'h00002864 : data <= 8'b00000000 ;
			15'h00002865 : data <= 8'b00000000 ;
			15'h00002866 : data <= 8'b00000000 ;
			15'h00002867 : data <= 8'b00000000 ;
			15'h00002868 : data <= 8'b00000000 ;
			15'h00002869 : data <= 8'b00000000 ;
			15'h0000286A : data <= 8'b00000000 ;
			15'h0000286B : data <= 8'b00000000 ;
			15'h0000286C : data <= 8'b00000000 ;
			15'h0000286D : data <= 8'b00000000 ;
			15'h0000286E : data <= 8'b00000000 ;
			15'h0000286F : data <= 8'b00000000 ;
			15'h00002870 : data <= 8'b00000000 ;
			15'h00002871 : data <= 8'b00000000 ;
			15'h00002872 : data <= 8'b00000000 ;
			15'h00002873 : data <= 8'b00000000 ;
			15'h00002874 : data <= 8'b00000000 ;
			15'h00002875 : data <= 8'b00000000 ;
			15'h00002876 : data <= 8'b00000000 ;
			15'h00002877 : data <= 8'b00000000 ;
			15'h00002878 : data <= 8'b00000000 ;
			15'h00002879 : data <= 8'b00000000 ;
			15'h0000287A : data <= 8'b00000000 ;
			15'h0000287B : data <= 8'b00000000 ;
			15'h0000287C : data <= 8'b00000000 ;
			15'h0000287D : data <= 8'b00000000 ;
			15'h0000287E : data <= 8'b00000000 ;
			15'h0000287F : data <= 8'b00000000 ;
			15'h00002880 : data <= 8'b00000000 ;
			15'h00002881 : data <= 8'b00000000 ;
			15'h00002882 : data <= 8'b00000000 ;
			15'h00002883 : data <= 8'b00000000 ;
			15'h00002884 : data <= 8'b00000000 ;
			15'h00002885 : data <= 8'b00000000 ;
			15'h00002886 : data <= 8'b00000000 ;
			15'h00002887 : data <= 8'b00000000 ;
			15'h00002888 : data <= 8'b00000000 ;
			15'h00002889 : data <= 8'b00000000 ;
			15'h0000288A : data <= 8'b00000000 ;
			15'h0000288B : data <= 8'b00000000 ;
			15'h0000288C : data <= 8'b00000000 ;
			15'h0000288D : data <= 8'b00000000 ;
			15'h0000288E : data <= 8'b00000000 ;
			15'h0000288F : data <= 8'b00000000 ;
			15'h00002890 : data <= 8'b00000000 ;
			15'h00002891 : data <= 8'b00000000 ;
			15'h00002892 : data <= 8'b00000000 ;
			15'h00002893 : data <= 8'b00000000 ;
			15'h00002894 : data <= 8'b00000000 ;
			15'h00002895 : data <= 8'b00000000 ;
			15'h00002896 : data <= 8'b00000000 ;
			15'h00002897 : data <= 8'b00000000 ;
			15'h00002898 : data <= 8'b00000000 ;
			15'h00002899 : data <= 8'b00000000 ;
			15'h0000289A : data <= 8'b00000000 ;
			15'h0000289B : data <= 8'b00000000 ;
			15'h0000289C : data <= 8'b00000000 ;
			15'h0000289D : data <= 8'b00000000 ;
			15'h0000289E : data <= 8'b00000000 ;
			15'h0000289F : data <= 8'b00000000 ;
			15'h000028A0 : data <= 8'b00000000 ;
			15'h000028A1 : data <= 8'b00000000 ;
			15'h000028A2 : data <= 8'b00000000 ;
			15'h000028A3 : data <= 8'b00000000 ;
			15'h000028A4 : data <= 8'b00000000 ;
			15'h000028A5 : data <= 8'b00000000 ;
			15'h000028A6 : data <= 8'b00000000 ;
			15'h000028A7 : data <= 8'b00000000 ;
			15'h000028A8 : data <= 8'b00000000 ;
			15'h000028A9 : data <= 8'b00000000 ;
			15'h000028AA : data <= 8'b00000000 ;
			15'h000028AB : data <= 8'b00000000 ;
			15'h000028AC : data <= 8'b00000000 ;
			15'h000028AD : data <= 8'b00000000 ;
			15'h000028AE : data <= 8'b00000000 ;
			15'h000028AF : data <= 8'b00000000 ;
			15'h000028B0 : data <= 8'b00000000 ;
			15'h000028B1 : data <= 8'b00000000 ;
			15'h000028B2 : data <= 8'b00000000 ;
			15'h000028B3 : data <= 8'b00000000 ;
			15'h000028B4 : data <= 8'b00000000 ;
			15'h000028B5 : data <= 8'b00000000 ;
			15'h000028B6 : data <= 8'b00000000 ;
			15'h000028B7 : data <= 8'b00000000 ;
			15'h000028B8 : data <= 8'b00000000 ;
			15'h000028B9 : data <= 8'b00000000 ;
			15'h000028BA : data <= 8'b00000000 ;
			15'h000028BB : data <= 8'b00000000 ;
			15'h000028BC : data <= 8'b00000000 ;
			15'h000028BD : data <= 8'b00000000 ;
			15'h000028BE : data <= 8'b00000000 ;
			15'h000028BF : data <= 8'b00000000 ;
			15'h000028C0 : data <= 8'b00000000 ;
			15'h000028C1 : data <= 8'b00000000 ;
			15'h000028C2 : data <= 8'b00000000 ;
			15'h000028C3 : data <= 8'b00000000 ;
			15'h000028C4 : data <= 8'b00000000 ;
			15'h000028C5 : data <= 8'b00000000 ;
			15'h000028C6 : data <= 8'b00000000 ;
			15'h000028C7 : data <= 8'b00000000 ;
			15'h000028C8 : data <= 8'b00000000 ;
			15'h000028C9 : data <= 8'b00000000 ;
			15'h000028CA : data <= 8'b00000000 ;
			15'h000028CB : data <= 8'b00000000 ;
			15'h000028CC : data <= 8'b00000000 ;
			15'h000028CD : data <= 8'b00000000 ;
			15'h000028CE : data <= 8'b00000000 ;
			15'h000028CF : data <= 8'b00000000 ;
			15'h000028D0 : data <= 8'b00000000 ;
			15'h000028D1 : data <= 8'b00000000 ;
			15'h000028D2 : data <= 8'b00000000 ;
			15'h000028D3 : data <= 8'b00000000 ;
			15'h000028D4 : data <= 8'b00000000 ;
			15'h000028D5 : data <= 8'b00000000 ;
			15'h000028D6 : data <= 8'b00000000 ;
			15'h000028D7 : data <= 8'b00000000 ;
			15'h000028D8 : data <= 8'b00000000 ;
			15'h000028D9 : data <= 8'b00000000 ;
			15'h000028DA : data <= 8'b00000000 ;
			15'h000028DB : data <= 8'b00000000 ;
			15'h000028DC : data <= 8'b00000000 ;
			15'h000028DD : data <= 8'b00000000 ;
			15'h000028DE : data <= 8'b00000000 ;
			15'h000028DF : data <= 8'b00000000 ;
			15'h000028E0 : data <= 8'b00000000 ;
			15'h000028E1 : data <= 8'b00000000 ;
			15'h000028E2 : data <= 8'b00000000 ;
			15'h000028E3 : data <= 8'b00000000 ;
			15'h000028E4 : data <= 8'b00000000 ;
			15'h000028E5 : data <= 8'b00000000 ;
			15'h000028E6 : data <= 8'b00000000 ;
			15'h000028E7 : data <= 8'b00000000 ;
			15'h000028E8 : data <= 8'b00000000 ;
			15'h000028E9 : data <= 8'b00000000 ;
			15'h000028EA : data <= 8'b00000000 ;
			15'h000028EB : data <= 8'b00000000 ;
			15'h000028EC : data <= 8'b00000000 ;
			15'h000028ED : data <= 8'b00000000 ;
			15'h000028EE : data <= 8'b00000000 ;
			15'h000028EF : data <= 8'b00000000 ;
			15'h000028F0 : data <= 8'b00000000 ;
			15'h000028F1 : data <= 8'b00000000 ;
			15'h000028F2 : data <= 8'b00000000 ;
			15'h000028F3 : data <= 8'b00000000 ;
			15'h000028F4 : data <= 8'b00000000 ;
			15'h000028F5 : data <= 8'b00000000 ;
			15'h000028F6 : data <= 8'b00000000 ;
			15'h000028F7 : data <= 8'b00000000 ;
			15'h000028F8 : data <= 8'b00000000 ;
			15'h000028F9 : data <= 8'b00000000 ;
			15'h000028FA : data <= 8'b00000000 ;
			15'h000028FB : data <= 8'b00000000 ;
			15'h000028FC : data <= 8'b00000000 ;
			15'h000028FD : data <= 8'b00000000 ;
			15'h000028FE : data <= 8'b00000000 ;
			15'h000028FF : data <= 8'b00000000 ;
			15'h00002900 : data <= 8'b00000000 ;
			15'h00002901 : data <= 8'b00000000 ;
			15'h00002902 : data <= 8'b00000000 ;
			15'h00002903 : data <= 8'b00000000 ;
			15'h00002904 : data <= 8'b00000000 ;
			15'h00002905 : data <= 8'b00000000 ;
			15'h00002906 : data <= 8'b00000000 ;
			15'h00002907 : data <= 8'b00000000 ;
			15'h00002908 : data <= 8'b00000000 ;
			15'h00002909 : data <= 8'b00000000 ;
			15'h0000290A : data <= 8'b00000000 ;
			15'h0000290B : data <= 8'b00000000 ;
			15'h0000290C : data <= 8'b00000000 ;
			15'h0000290D : data <= 8'b00000000 ;
			15'h0000290E : data <= 8'b00000000 ;
			15'h0000290F : data <= 8'b00000000 ;
			15'h00002910 : data <= 8'b00000000 ;
			15'h00002911 : data <= 8'b00000000 ;
			15'h00002912 : data <= 8'b00000000 ;
			15'h00002913 : data <= 8'b00000000 ;
			15'h00002914 : data <= 8'b00000000 ;
			15'h00002915 : data <= 8'b00000000 ;
			15'h00002916 : data <= 8'b00000000 ;
			15'h00002917 : data <= 8'b00000000 ;
			15'h00002918 : data <= 8'b00000000 ;
			15'h00002919 : data <= 8'b00000000 ;
			15'h0000291A : data <= 8'b00000000 ;
			15'h0000291B : data <= 8'b00000000 ;
			15'h0000291C : data <= 8'b00000000 ;
			15'h0000291D : data <= 8'b00000000 ;
			15'h0000291E : data <= 8'b00000000 ;
			15'h0000291F : data <= 8'b00000000 ;
			15'h00002920 : data <= 8'b00000000 ;
			15'h00002921 : data <= 8'b00000000 ;
			15'h00002922 : data <= 8'b00000000 ;
			15'h00002923 : data <= 8'b00000000 ;
			15'h00002924 : data <= 8'b00000000 ;
			15'h00002925 : data <= 8'b00000000 ;
			15'h00002926 : data <= 8'b00000000 ;
			15'h00002927 : data <= 8'b00000000 ;
			15'h00002928 : data <= 8'b00000000 ;
			15'h00002929 : data <= 8'b00000000 ;
			15'h0000292A : data <= 8'b00000000 ;
			15'h0000292B : data <= 8'b00000000 ;
			15'h0000292C : data <= 8'b00000000 ;
			15'h0000292D : data <= 8'b00000000 ;
			15'h0000292E : data <= 8'b00000000 ;
			15'h0000292F : data <= 8'b00000000 ;
			15'h00002930 : data <= 8'b00000000 ;
			15'h00002931 : data <= 8'b00000000 ;
			15'h00002932 : data <= 8'b00000000 ;
			15'h00002933 : data <= 8'b00000000 ;
			15'h00002934 : data <= 8'b00000000 ;
			15'h00002935 : data <= 8'b00000000 ;
			15'h00002936 : data <= 8'b00000000 ;
			15'h00002937 : data <= 8'b00000000 ;
			15'h00002938 : data <= 8'b00000000 ;
			15'h00002939 : data <= 8'b00000000 ;
			15'h0000293A : data <= 8'b00000000 ;
			15'h0000293B : data <= 8'b00000000 ;
			15'h0000293C : data <= 8'b00000000 ;
			15'h0000293D : data <= 8'b00000000 ;
			15'h0000293E : data <= 8'b00000000 ;
			15'h0000293F : data <= 8'b00000000 ;
			15'h00002940 : data <= 8'b00000000 ;
			15'h00002941 : data <= 8'b00000000 ;
			15'h00002942 : data <= 8'b00000000 ;
			15'h00002943 : data <= 8'b00000000 ;
			15'h00002944 : data <= 8'b00000000 ;
			15'h00002945 : data <= 8'b00000000 ;
			15'h00002946 : data <= 8'b00000000 ;
			15'h00002947 : data <= 8'b00000000 ;
			15'h00002948 : data <= 8'b00000000 ;
			15'h00002949 : data <= 8'b00000000 ;
			15'h0000294A : data <= 8'b00000000 ;
			15'h0000294B : data <= 8'b00000000 ;
			15'h0000294C : data <= 8'b00000000 ;
			15'h0000294D : data <= 8'b00000000 ;
			15'h0000294E : data <= 8'b00000000 ;
			15'h0000294F : data <= 8'b00000000 ;
			15'h00002950 : data <= 8'b00000000 ;
			15'h00002951 : data <= 8'b00000000 ;
			15'h00002952 : data <= 8'b00000000 ;
			15'h00002953 : data <= 8'b00000000 ;
			15'h00002954 : data <= 8'b00000000 ;
			15'h00002955 : data <= 8'b00000000 ;
			15'h00002956 : data <= 8'b00000000 ;
			15'h00002957 : data <= 8'b00000000 ;
			15'h00002958 : data <= 8'b00000000 ;
			15'h00002959 : data <= 8'b00000000 ;
			15'h0000295A : data <= 8'b00000000 ;
			15'h0000295B : data <= 8'b00000000 ;
			15'h0000295C : data <= 8'b00000000 ;
			15'h0000295D : data <= 8'b00000000 ;
			15'h0000295E : data <= 8'b00000000 ;
			15'h0000295F : data <= 8'b00000000 ;
			15'h00002960 : data <= 8'b00000000 ;
			15'h00002961 : data <= 8'b00000000 ;
			15'h00002962 : data <= 8'b00000000 ;
			15'h00002963 : data <= 8'b00000000 ;
			15'h00002964 : data <= 8'b00000000 ;
			15'h00002965 : data <= 8'b00000000 ;
			15'h00002966 : data <= 8'b00000000 ;
			15'h00002967 : data <= 8'b00000000 ;
			15'h00002968 : data <= 8'b00000000 ;
			15'h00002969 : data <= 8'b00000000 ;
			15'h0000296A : data <= 8'b00000000 ;
			15'h0000296B : data <= 8'b00000000 ;
			15'h0000296C : data <= 8'b00000000 ;
			15'h0000296D : data <= 8'b00000000 ;
			15'h0000296E : data <= 8'b00000000 ;
			15'h0000296F : data <= 8'b00000000 ;
			15'h00002970 : data <= 8'b00000000 ;
			15'h00002971 : data <= 8'b00000000 ;
			15'h00002972 : data <= 8'b00000000 ;
			15'h00002973 : data <= 8'b00000000 ;
			15'h00002974 : data <= 8'b00000000 ;
			15'h00002975 : data <= 8'b00000000 ;
			15'h00002976 : data <= 8'b00000000 ;
			15'h00002977 : data <= 8'b00000000 ;
			15'h00002978 : data <= 8'b00000000 ;
			15'h00002979 : data <= 8'b00000000 ;
			15'h0000297A : data <= 8'b00000000 ;
			15'h0000297B : data <= 8'b00000000 ;
			15'h0000297C : data <= 8'b00000000 ;
			15'h0000297D : data <= 8'b00000000 ;
			15'h0000297E : data <= 8'b00000000 ;
			15'h0000297F : data <= 8'b00000000 ;
			15'h00002980 : data <= 8'b00000000 ;
			15'h00002981 : data <= 8'b00000000 ;
			15'h00002982 : data <= 8'b00000000 ;
			15'h00002983 : data <= 8'b00000000 ;
			15'h00002984 : data <= 8'b00000000 ;
			15'h00002985 : data <= 8'b00000000 ;
			15'h00002986 : data <= 8'b00000000 ;
			15'h00002987 : data <= 8'b00000000 ;
			15'h00002988 : data <= 8'b00000000 ;
			15'h00002989 : data <= 8'b00000000 ;
			15'h0000298A : data <= 8'b00000000 ;
			15'h0000298B : data <= 8'b00000000 ;
			15'h0000298C : data <= 8'b00000000 ;
			15'h0000298D : data <= 8'b00000000 ;
			15'h0000298E : data <= 8'b00000000 ;
			15'h0000298F : data <= 8'b00000000 ;
			15'h00002990 : data <= 8'b00000000 ;
			15'h00002991 : data <= 8'b00000000 ;
			15'h00002992 : data <= 8'b00000000 ;
			15'h00002993 : data <= 8'b00000000 ;
			15'h00002994 : data <= 8'b00000000 ;
			15'h00002995 : data <= 8'b00000000 ;
			15'h00002996 : data <= 8'b00000000 ;
			15'h00002997 : data <= 8'b00000000 ;
			15'h00002998 : data <= 8'b00000000 ;
			15'h00002999 : data <= 8'b00000000 ;
			15'h0000299A : data <= 8'b00000000 ;
			15'h0000299B : data <= 8'b00000000 ;
			15'h0000299C : data <= 8'b00000000 ;
			15'h0000299D : data <= 8'b00000000 ;
			15'h0000299E : data <= 8'b00000000 ;
			15'h0000299F : data <= 8'b00000000 ;
			15'h000029A0 : data <= 8'b00000000 ;
			15'h000029A1 : data <= 8'b00000000 ;
			15'h000029A2 : data <= 8'b00000000 ;
			15'h000029A3 : data <= 8'b00000000 ;
			15'h000029A4 : data <= 8'b00000000 ;
			15'h000029A5 : data <= 8'b00000000 ;
			15'h000029A6 : data <= 8'b00000000 ;
			15'h000029A7 : data <= 8'b00000000 ;
			15'h000029A8 : data <= 8'b00000000 ;
			15'h000029A9 : data <= 8'b00000000 ;
			15'h000029AA : data <= 8'b00000000 ;
			15'h000029AB : data <= 8'b00000000 ;
			15'h000029AC : data <= 8'b00000000 ;
			15'h000029AD : data <= 8'b00000000 ;
			15'h000029AE : data <= 8'b00000000 ;
			15'h000029AF : data <= 8'b00000000 ;
			15'h000029B0 : data <= 8'b00000000 ;
			15'h000029B1 : data <= 8'b00000000 ;
			15'h000029B2 : data <= 8'b00000000 ;
			15'h000029B3 : data <= 8'b00000000 ;
			15'h000029B4 : data <= 8'b00000000 ;
			15'h000029B5 : data <= 8'b00000000 ;
			15'h000029B6 : data <= 8'b00000000 ;
			15'h000029B7 : data <= 8'b00000000 ;
			15'h000029B8 : data <= 8'b00000000 ;
			15'h000029B9 : data <= 8'b00000000 ;
			15'h000029BA : data <= 8'b00000000 ;
			15'h000029BB : data <= 8'b00000000 ;
			15'h000029BC : data <= 8'b00000000 ;
			15'h000029BD : data <= 8'b00000000 ;
			15'h000029BE : data <= 8'b00000000 ;
			15'h000029BF : data <= 8'b00000000 ;
			15'h000029C0 : data <= 8'b00000000 ;
			15'h000029C1 : data <= 8'b00000000 ;
			15'h000029C2 : data <= 8'b00000000 ;
			15'h000029C3 : data <= 8'b00000000 ;
			15'h000029C4 : data <= 8'b00000000 ;
			15'h000029C5 : data <= 8'b00000000 ;
			15'h000029C6 : data <= 8'b00000000 ;
			15'h000029C7 : data <= 8'b00000000 ;
			15'h000029C8 : data <= 8'b00000000 ;
			15'h000029C9 : data <= 8'b00000000 ;
			15'h000029CA : data <= 8'b00000000 ;
			15'h000029CB : data <= 8'b00000000 ;
			15'h000029CC : data <= 8'b00000000 ;
			15'h000029CD : data <= 8'b00000000 ;
			15'h000029CE : data <= 8'b00000000 ;
			15'h000029CF : data <= 8'b00000000 ;
			15'h000029D0 : data <= 8'b00000000 ;
			15'h000029D1 : data <= 8'b00000000 ;
			15'h000029D2 : data <= 8'b00000000 ;
			15'h000029D3 : data <= 8'b00000000 ;
			15'h000029D4 : data <= 8'b00000000 ;
			15'h000029D5 : data <= 8'b00000000 ;
			15'h000029D6 : data <= 8'b00000000 ;
			15'h000029D7 : data <= 8'b00000000 ;
			15'h000029D8 : data <= 8'b00000000 ;
			15'h000029D9 : data <= 8'b00000000 ;
			15'h000029DA : data <= 8'b00000000 ;
			15'h000029DB : data <= 8'b00000000 ;
			15'h000029DC : data <= 8'b00000000 ;
			15'h000029DD : data <= 8'b00000000 ;
			15'h000029DE : data <= 8'b00000000 ;
			15'h000029DF : data <= 8'b00000000 ;
			15'h000029E0 : data <= 8'b00000000 ;
			15'h000029E1 : data <= 8'b00000000 ;
			15'h000029E2 : data <= 8'b00000000 ;
			15'h000029E3 : data <= 8'b00000000 ;
			15'h000029E4 : data <= 8'b00000000 ;
			15'h000029E5 : data <= 8'b00000000 ;
			15'h000029E6 : data <= 8'b00000000 ;
			15'h000029E7 : data <= 8'b00000000 ;
			15'h000029E8 : data <= 8'b00000000 ;
			15'h000029E9 : data <= 8'b00000000 ;
			15'h000029EA : data <= 8'b00000000 ;
			15'h000029EB : data <= 8'b00000000 ;
			15'h000029EC : data <= 8'b00000000 ;
			15'h000029ED : data <= 8'b00000000 ;
			15'h000029EE : data <= 8'b00000000 ;
			15'h000029EF : data <= 8'b00000000 ;
			15'h000029F0 : data <= 8'b00000000 ;
			15'h000029F1 : data <= 8'b00000000 ;
			15'h000029F2 : data <= 8'b00000000 ;
			15'h000029F3 : data <= 8'b00000000 ;
			15'h000029F4 : data <= 8'b00000000 ;
			15'h000029F5 : data <= 8'b00000000 ;
			15'h000029F6 : data <= 8'b00000000 ;
			15'h000029F7 : data <= 8'b00000000 ;
			15'h000029F8 : data <= 8'b00000000 ;
			15'h000029F9 : data <= 8'b00000000 ;
			15'h000029FA : data <= 8'b00000000 ;
			15'h000029FB : data <= 8'b00000000 ;
			15'h000029FC : data <= 8'b00000000 ;
			15'h000029FD : data <= 8'b00000000 ;
			15'h000029FE : data <= 8'b00000000 ;
			15'h000029FF : data <= 8'b00000000 ;
			15'h00002A00 : data <= 8'b00000000 ;
			15'h00002A01 : data <= 8'b00000000 ;
			15'h00002A02 : data <= 8'b00000000 ;
			15'h00002A03 : data <= 8'b00000000 ;
			15'h00002A04 : data <= 8'b00000000 ;
			15'h00002A05 : data <= 8'b00000000 ;
			15'h00002A06 : data <= 8'b00000000 ;
			15'h00002A07 : data <= 8'b00000000 ;
			15'h00002A08 : data <= 8'b00000000 ;
			15'h00002A09 : data <= 8'b00000000 ;
			15'h00002A0A : data <= 8'b00000000 ;
			15'h00002A0B : data <= 8'b00000000 ;
			15'h00002A0C : data <= 8'b00000000 ;
			15'h00002A0D : data <= 8'b00000000 ;
			15'h00002A0E : data <= 8'b00000000 ;
			15'h00002A0F : data <= 8'b00000000 ;
			15'h00002A10 : data <= 8'b00000000 ;
			15'h00002A11 : data <= 8'b00000000 ;
			15'h00002A12 : data <= 8'b00000000 ;
			15'h00002A13 : data <= 8'b00000000 ;
			15'h00002A14 : data <= 8'b00000000 ;
			15'h00002A15 : data <= 8'b00000000 ;
			15'h00002A16 : data <= 8'b00000000 ;
			15'h00002A17 : data <= 8'b00000000 ;
			15'h00002A18 : data <= 8'b00000000 ;
			15'h00002A19 : data <= 8'b00000000 ;
			15'h00002A1A : data <= 8'b00000000 ;
			15'h00002A1B : data <= 8'b00000000 ;
			15'h00002A1C : data <= 8'b00000000 ;
			15'h00002A1D : data <= 8'b00000000 ;
			15'h00002A1E : data <= 8'b00000000 ;
			15'h00002A1F : data <= 8'b00000000 ;
			15'h00002A20 : data <= 8'b00000000 ;
			15'h00002A21 : data <= 8'b00000000 ;
			15'h00002A22 : data <= 8'b00000000 ;
			15'h00002A23 : data <= 8'b00000000 ;
			15'h00002A24 : data <= 8'b00000000 ;
			15'h00002A25 : data <= 8'b00000000 ;
			15'h00002A26 : data <= 8'b00000000 ;
			15'h00002A27 : data <= 8'b00000000 ;
			15'h00002A28 : data <= 8'b00000000 ;
			15'h00002A29 : data <= 8'b00000000 ;
			15'h00002A2A : data <= 8'b00000000 ;
			15'h00002A2B : data <= 8'b00000000 ;
			15'h00002A2C : data <= 8'b00000000 ;
			15'h00002A2D : data <= 8'b00000000 ;
			15'h00002A2E : data <= 8'b00000000 ;
			15'h00002A2F : data <= 8'b00000000 ;
			15'h00002A30 : data <= 8'b00000000 ;
			15'h00002A31 : data <= 8'b00000000 ;
			15'h00002A32 : data <= 8'b00000000 ;
			15'h00002A33 : data <= 8'b00000000 ;
			15'h00002A34 : data <= 8'b00000000 ;
			15'h00002A35 : data <= 8'b00000000 ;
			15'h00002A36 : data <= 8'b00000000 ;
			15'h00002A37 : data <= 8'b00000000 ;
			15'h00002A38 : data <= 8'b00000000 ;
			15'h00002A39 : data <= 8'b00000000 ;
			15'h00002A3A : data <= 8'b00000000 ;
			15'h00002A3B : data <= 8'b00000000 ;
			15'h00002A3C : data <= 8'b00000000 ;
			15'h00002A3D : data <= 8'b00000000 ;
			15'h00002A3E : data <= 8'b00000000 ;
			15'h00002A3F : data <= 8'b00000000 ;
			15'h00002A40 : data <= 8'b00000000 ;
			15'h00002A41 : data <= 8'b00000000 ;
			15'h00002A42 : data <= 8'b00000000 ;
			15'h00002A43 : data <= 8'b00000000 ;
			15'h00002A44 : data <= 8'b00000000 ;
			15'h00002A45 : data <= 8'b00000000 ;
			15'h00002A46 : data <= 8'b00000000 ;
			15'h00002A47 : data <= 8'b00000000 ;
			15'h00002A48 : data <= 8'b00000000 ;
			15'h00002A49 : data <= 8'b00000000 ;
			15'h00002A4A : data <= 8'b00000000 ;
			15'h00002A4B : data <= 8'b00000000 ;
			15'h00002A4C : data <= 8'b00000000 ;
			15'h00002A4D : data <= 8'b00000000 ;
			15'h00002A4E : data <= 8'b00000000 ;
			15'h00002A4F : data <= 8'b00000000 ;
			15'h00002A50 : data <= 8'b00000000 ;
			15'h00002A51 : data <= 8'b00000000 ;
			15'h00002A52 : data <= 8'b00000000 ;
			15'h00002A53 : data <= 8'b00000000 ;
			15'h00002A54 : data <= 8'b00000000 ;
			15'h00002A55 : data <= 8'b00000000 ;
			15'h00002A56 : data <= 8'b00000000 ;
			15'h00002A57 : data <= 8'b00000000 ;
			15'h00002A58 : data <= 8'b00000000 ;
			15'h00002A59 : data <= 8'b00000000 ;
			15'h00002A5A : data <= 8'b00000000 ;
			15'h00002A5B : data <= 8'b00000000 ;
			15'h00002A5C : data <= 8'b00000000 ;
			15'h00002A5D : data <= 8'b00000000 ;
			15'h00002A5E : data <= 8'b00000000 ;
			15'h00002A5F : data <= 8'b00000000 ;
			15'h00002A60 : data <= 8'b00000000 ;
			15'h00002A61 : data <= 8'b00000000 ;
			15'h00002A62 : data <= 8'b00000000 ;
			15'h00002A63 : data <= 8'b00000000 ;
			15'h00002A64 : data <= 8'b00000000 ;
			15'h00002A65 : data <= 8'b00000000 ;
			15'h00002A66 : data <= 8'b00000000 ;
			15'h00002A67 : data <= 8'b00000000 ;
			15'h00002A68 : data <= 8'b00000000 ;
			15'h00002A69 : data <= 8'b00000000 ;
			15'h00002A6A : data <= 8'b00000000 ;
			15'h00002A6B : data <= 8'b00000000 ;
			15'h00002A6C : data <= 8'b00000000 ;
			15'h00002A6D : data <= 8'b00000000 ;
			15'h00002A6E : data <= 8'b00000000 ;
			15'h00002A6F : data <= 8'b00000000 ;
			15'h00002A70 : data <= 8'b00000000 ;
			15'h00002A71 : data <= 8'b00000000 ;
			15'h00002A72 : data <= 8'b00000000 ;
			15'h00002A73 : data <= 8'b00000000 ;
			15'h00002A74 : data <= 8'b00000000 ;
			15'h00002A75 : data <= 8'b00000000 ;
			15'h00002A76 : data <= 8'b00000000 ;
			15'h00002A77 : data <= 8'b00000000 ;
			15'h00002A78 : data <= 8'b00000000 ;
			15'h00002A79 : data <= 8'b00000000 ;
			15'h00002A7A : data <= 8'b00000000 ;
			15'h00002A7B : data <= 8'b00000000 ;
			15'h00002A7C : data <= 8'b00000000 ;
			15'h00002A7D : data <= 8'b00000000 ;
			15'h00002A7E : data <= 8'b00000000 ;
			15'h00002A7F : data <= 8'b00000000 ;
			15'h00002A80 : data <= 8'b00000000 ;
			15'h00002A81 : data <= 8'b00000000 ;
			15'h00002A82 : data <= 8'b00000000 ;
			15'h00002A83 : data <= 8'b00000000 ;
			15'h00002A84 : data <= 8'b00000000 ;
			15'h00002A85 : data <= 8'b00000000 ;
			15'h00002A86 : data <= 8'b00000000 ;
			15'h00002A87 : data <= 8'b00000000 ;
			15'h00002A88 : data <= 8'b00000000 ;
			15'h00002A89 : data <= 8'b00000000 ;
			15'h00002A8A : data <= 8'b00000000 ;
			15'h00002A8B : data <= 8'b00000000 ;
			15'h00002A8C : data <= 8'b00000000 ;
			15'h00002A8D : data <= 8'b00000000 ;
			15'h00002A8E : data <= 8'b00000000 ;
			15'h00002A8F : data <= 8'b00000000 ;
			15'h00002A90 : data <= 8'b00000000 ;
			15'h00002A91 : data <= 8'b00000000 ;
			15'h00002A92 : data <= 8'b00000000 ;
			15'h00002A93 : data <= 8'b00000000 ;
			15'h00002A94 : data <= 8'b00000000 ;
			15'h00002A95 : data <= 8'b00000000 ;
			15'h00002A96 : data <= 8'b00000000 ;
			15'h00002A97 : data <= 8'b00000000 ;
			15'h00002A98 : data <= 8'b00000000 ;
			15'h00002A99 : data <= 8'b00000000 ;
			15'h00002A9A : data <= 8'b00000000 ;
			15'h00002A9B : data <= 8'b00000000 ;
			15'h00002A9C : data <= 8'b00000000 ;
			15'h00002A9D : data <= 8'b00000000 ;
			15'h00002A9E : data <= 8'b00000000 ;
			15'h00002A9F : data <= 8'b00000000 ;
			15'h00002AA0 : data <= 8'b00000000 ;
			15'h00002AA1 : data <= 8'b00000000 ;
			15'h00002AA2 : data <= 8'b00000000 ;
			15'h00002AA3 : data <= 8'b00000000 ;
			15'h00002AA4 : data <= 8'b00000000 ;
			15'h00002AA5 : data <= 8'b00000000 ;
			15'h00002AA6 : data <= 8'b00000000 ;
			15'h00002AA7 : data <= 8'b00000000 ;
			15'h00002AA8 : data <= 8'b00000000 ;
			15'h00002AA9 : data <= 8'b00000000 ;
			15'h00002AAA : data <= 8'b00000000 ;
			15'h00002AAB : data <= 8'b00000000 ;
			15'h00002AAC : data <= 8'b00000000 ;
			15'h00002AAD : data <= 8'b00000000 ;
			15'h00002AAE : data <= 8'b00000000 ;
			15'h00002AAF : data <= 8'b00000000 ;
			15'h00002AB0 : data <= 8'b00000000 ;
			15'h00002AB1 : data <= 8'b00000000 ;
			15'h00002AB2 : data <= 8'b00000000 ;
			15'h00002AB3 : data <= 8'b00000000 ;
			15'h00002AB4 : data <= 8'b00000000 ;
			15'h00002AB5 : data <= 8'b00000000 ;
			15'h00002AB6 : data <= 8'b00000000 ;
			15'h00002AB7 : data <= 8'b00000000 ;
			15'h00002AB8 : data <= 8'b00000000 ;
			15'h00002AB9 : data <= 8'b00000000 ;
			15'h00002ABA : data <= 8'b00000000 ;
			15'h00002ABB : data <= 8'b00000000 ;
			15'h00002ABC : data <= 8'b00000000 ;
			15'h00002ABD : data <= 8'b00000000 ;
			15'h00002ABE : data <= 8'b00000000 ;
			15'h00002ABF : data <= 8'b00000000 ;
			15'h00002AC0 : data <= 8'b00000000 ;
			15'h00002AC1 : data <= 8'b00000000 ;
			15'h00002AC2 : data <= 8'b00000000 ;
			15'h00002AC3 : data <= 8'b00000000 ;
			15'h00002AC4 : data <= 8'b00000000 ;
			15'h00002AC5 : data <= 8'b00000000 ;
			15'h00002AC6 : data <= 8'b00000000 ;
			15'h00002AC7 : data <= 8'b00000000 ;
			15'h00002AC8 : data <= 8'b00000000 ;
			15'h00002AC9 : data <= 8'b00000000 ;
			15'h00002ACA : data <= 8'b00000000 ;
			15'h00002ACB : data <= 8'b00000000 ;
			15'h00002ACC : data <= 8'b00000000 ;
			15'h00002ACD : data <= 8'b00000000 ;
			15'h00002ACE : data <= 8'b00000000 ;
			15'h00002ACF : data <= 8'b00000000 ;
			15'h00002AD0 : data <= 8'b00000000 ;
			15'h00002AD1 : data <= 8'b00000000 ;
			15'h00002AD2 : data <= 8'b00000000 ;
			15'h00002AD3 : data <= 8'b00000000 ;
			15'h00002AD4 : data <= 8'b00000000 ;
			15'h00002AD5 : data <= 8'b00000000 ;
			15'h00002AD6 : data <= 8'b00000000 ;
			15'h00002AD7 : data <= 8'b00000000 ;
			15'h00002AD8 : data <= 8'b00000000 ;
			15'h00002AD9 : data <= 8'b00000000 ;
			15'h00002ADA : data <= 8'b00000000 ;
			15'h00002ADB : data <= 8'b00000000 ;
			15'h00002ADC : data <= 8'b00000000 ;
			15'h00002ADD : data <= 8'b00000000 ;
			15'h00002ADE : data <= 8'b00000000 ;
			15'h00002ADF : data <= 8'b00000000 ;
			15'h00002AE0 : data <= 8'b00000000 ;
			15'h00002AE1 : data <= 8'b00000000 ;
			15'h00002AE2 : data <= 8'b00000000 ;
			15'h00002AE3 : data <= 8'b00000000 ;
			15'h00002AE4 : data <= 8'b00000000 ;
			15'h00002AE5 : data <= 8'b00000000 ;
			15'h00002AE6 : data <= 8'b00000000 ;
			15'h00002AE7 : data <= 8'b00000000 ;
			15'h00002AE8 : data <= 8'b00000000 ;
			15'h00002AE9 : data <= 8'b00000000 ;
			15'h00002AEA : data <= 8'b00000000 ;
			15'h00002AEB : data <= 8'b00000000 ;
			15'h00002AEC : data <= 8'b00000000 ;
			15'h00002AED : data <= 8'b00000000 ;
			15'h00002AEE : data <= 8'b00000000 ;
			15'h00002AEF : data <= 8'b00000000 ;
			15'h00002AF0 : data <= 8'b00000000 ;
			15'h00002AF1 : data <= 8'b00000000 ;
			15'h00002AF2 : data <= 8'b00000000 ;
			15'h00002AF3 : data <= 8'b00000000 ;
			15'h00002AF4 : data <= 8'b00000000 ;
			15'h00002AF5 : data <= 8'b00000000 ;
			15'h00002AF6 : data <= 8'b00000000 ;
			15'h00002AF7 : data <= 8'b00000000 ;
			15'h00002AF8 : data <= 8'b00000000 ;
			15'h00002AF9 : data <= 8'b00000000 ;
			15'h00002AFA : data <= 8'b00000000 ;
			15'h00002AFB : data <= 8'b00000000 ;
			15'h00002AFC : data <= 8'b00000000 ;
			15'h00002AFD : data <= 8'b00000000 ;
			15'h00002AFE : data <= 8'b00000000 ;
			15'h00002AFF : data <= 8'b00000000 ;
			15'h00002B00 : data <= 8'b00000000 ;
			15'h00002B01 : data <= 8'b00000000 ;
			15'h00002B02 : data <= 8'b00000000 ;
			15'h00002B03 : data <= 8'b00000000 ;
			15'h00002B04 : data <= 8'b00000000 ;
			15'h00002B05 : data <= 8'b00000000 ;
			15'h00002B06 : data <= 8'b00000000 ;
			15'h00002B07 : data <= 8'b00000000 ;
			15'h00002B08 : data <= 8'b00000000 ;
			15'h00002B09 : data <= 8'b00000000 ;
			15'h00002B0A : data <= 8'b00000000 ;
			15'h00002B0B : data <= 8'b00000000 ;
			15'h00002B0C : data <= 8'b00000000 ;
			15'h00002B0D : data <= 8'b00000000 ;
			15'h00002B0E : data <= 8'b00000000 ;
			15'h00002B0F : data <= 8'b00000000 ;
			15'h00002B10 : data <= 8'b00000000 ;
			15'h00002B11 : data <= 8'b00000000 ;
			15'h00002B12 : data <= 8'b00000000 ;
			15'h00002B13 : data <= 8'b00000000 ;
			15'h00002B14 : data <= 8'b00000000 ;
			15'h00002B15 : data <= 8'b00000000 ;
			15'h00002B16 : data <= 8'b00000000 ;
			15'h00002B17 : data <= 8'b00000000 ;
			15'h00002B18 : data <= 8'b00000000 ;
			15'h00002B19 : data <= 8'b00000000 ;
			15'h00002B1A : data <= 8'b00000000 ;
			15'h00002B1B : data <= 8'b00000000 ;
			15'h00002B1C : data <= 8'b00000000 ;
			15'h00002B1D : data <= 8'b00000000 ;
			15'h00002B1E : data <= 8'b00000000 ;
			15'h00002B1F : data <= 8'b00000000 ;
			15'h00002B20 : data <= 8'b00000000 ;
			15'h00002B21 : data <= 8'b00000000 ;
			15'h00002B22 : data <= 8'b00000000 ;
			15'h00002B23 : data <= 8'b00000000 ;
			15'h00002B24 : data <= 8'b00000000 ;
			15'h00002B25 : data <= 8'b00000000 ;
			15'h00002B26 : data <= 8'b00000000 ;
			15'h00002B27 : data <= 8'b00000000 ;
			15'h00002B28 : data <= 8'b00000000 ;
			15'h00002B29 : data <= 8'b00000000 ;
			15'h00002B2A : data <= 8'b00000000 ;
			15'h00002B2B : data <= 8'b00000000 ;
			15'h00002B2C : data <= 8'b00000000 ;
			15'h00002B2D : data <= 8'b00000000 ;
			15'h00002B2E : data <= 8'b00000000 ;
			15'h00002B2F : data <= 8'b00000000 ;
			15'h00002B30 : data <= 8'b00000000 ;
			15'h00002B31 : data <= 8'b00000000 ;
			15'h00002B32 : data <= 8'b00000000 ;
			15'h00002B33 : data <= 8'b00000000 ;
			15'h00002B34 : data <= 8'b00000000 ;
			15'h00002B35 : data <= 8'b00000000 ;
			15'h00002B36 : data <= 8'b00000000 ;
			15'h00002B37 : data <= 8'b00000000 ;
			15'h00002B38 : data <= 8'b00000000 ;
			15'h00002B39 : data <= 8'b00000000 ;
			15'h00002B3A : data <= 8'b00000000 ;
			15'h00002B3B : data <= 8'b00000000 ;
			15'h00002B3C : data <= 8'b00000000 ;
			15'h00002B3D : data <= 8'b00000000 ;
			15'h00002B3E : data <= 8'b00000000 ;
			15'h00002B3F : data <= 8'b00000000 ;
			15'h00002B40 : data <= 8'b00000000 ;
			15'h00002B41 : data <= 8'b00000000 ;
			15'h00002B42 : data <= 8'b00000000 ;
			15'h00002B43 : data <= 8'b00000000 ;
			15'h00002B44 : data <= 8'b00000000 ;
			15'h00002B45 : data <= 8'b00000000 ;
			15'h00002B46 : data <= 8'b00000000 ;
			15'h00002B47 : data <= 8'b00000000 ;
			15'h00002B48 : data <= 8'b00000000 ;
			15'h00002B49 : data <= 8'b00000000 ;
			15'h00002B4A : data <= 8'b00000000 ;
			15'h00002B4B : data <= 8'b00000000 ;
			15'h00002B4C : data <= 8'b00000000 ;
			15'h00002B4D : data <= 8'b00000000 ;
			15'h00002B4E : data <= 8'b00000000 ;
			15'h00002B4F : data <= 8'b00000000 ;
			15'h00002B50 : data <= 8'b00000000 ;
			15'h00002B51 : data <= 8'b00000000 ;
			15'h00002B52 : data <= 8'b00000000 ;
			15'h00002B53 : data <= 8'b00000000 ;
			15'h00002B54 : data <= 8'b00000000 ;
			15'h00002B55 : data <= 8'b00000000 ;
			15'h00002B56 : data <= 8'b00000000 ;
			15'h00002B57 : data <= 8'b00000000 ;
			15'h00002B58 : data <= 8'b00000000 ;
			15'h00002B59 : data <= 8'b00000000 ;
			15'h00002B5A : data <= 8'b00000000 ;
			15'h00002B5B : data <= 8'b00000000 ;
			15'h00002B5C : data <= 8'b00000000 ;
			15'h00002B5D : data <= 8'b00000000 ;
			15'h00002B5E : data <= 8'b00000000 ;
			15'h00002B5F : data <= 8'b00000000 ;
			15'h00002B60 : data <= 8'b00000000 ;
			15'h00002B61 : data <= 8'b00000000 ;
			15'h00002B62 : data <= 8'b00000000 ;
			15'h00002B63 : data <= 8'b00000000 ;
			15'h00002B64 : data <= 8'b00000000 ;
			15'h00002B65 : data <= 8'b00000000 ;
			15'h00002B66 : data <= 8'b00000000 ;
			15'h00002B67 : data <= 8'b00000000 ;
			15'h00002B68 : data <= 8'b00000000 ;
			15'h00002B69 : data <= 8'b00000000 ;
			15'h00002B6A : data <= 8'b00000000 ;
			15'h00002B6B : data <= 8'b00000000 ;
			15'h00002B6C : data <= 8'b00000000 ;
			15'h00002B6D : data <= 8'b00000000 ;
			15'h00002B6E : data <= 8'b00000000 ;
			15'h00002B6F : data <= 8'b00000000 ;
			15'h00002B70 : data <= 8'b00000000 ;
			15'h00002B71 : data <= 8'b00000000 ;
			15'h00002B72 : data <= 8'b00000000 ;
			15'h00002B73 : data <= 8'b00000000 ;
			15'h00002B74 : data <= 8'b00000000 ;
			15'h00002B75 : data <= 8'b00000000 ;
			15'h00002B76 : data <= 8'b00000000 ;
			15'h00002B77 : data <= 8'b00000000 ;
			15'h00002B78 : data <= 8'b00000000 ;
			15'h00002B79 : data <= 8'b00000000 ;
			15'h00002B7A : data <= 8'b00000000 ;
			15'h00002B7B : data <= 8'b00000000 ;
			15'h00002B7C : data <= 8'b00000000 ;
			15'h00002B7D : data <= 8'b00000000 ;
			15'h00002B7E : data <= 8'b00000000 ;
			15'h00002B7F : data <= 8'b00000000 ;
			15'h00002B80 : data <= 8'b00000000 ;
			15'h00002B81 : data <= 8'b00000000 ;
			15'h00002B82 : data <= 8'b00000000 ;
			15'h00002B83 : data <= 8'b00000000 ;
			15'h00002B84 : data <= 8'b00000000 ;
			15'h00002B85 : data <= 8'b00000000 ;
			15'h00002B86 : data <= 8'b00000000 ;
			15'h00002B87 : data <= 8'b00000000 ;
			15'h00002B88 : data <= 8'b00000000 ;
			15'h00002B89 : data <= 8'b00000000 ;
			15'h00002B8A : data <= 8'b00000000 ;
			15'h00002B8B : data <= 8'b00000000 ;
			15'h00002B8C : data <= 8'b00000000 ;
			15'h00002B8D : data <= 8'b00000000 ;
			15'h00002B8E : data <= 8'b00000000 ;
			15'h00002B8F : data <= 8'b00000000 ;
			15'h00002B90 : data <= 8'b00000000 ;
			15'h00002B91 : data <= 8'b00000000 ;
			15'h00002B92 : data <= 8'b00000000 ;
			15'h00002B93 : data <= 8'b00000000 ;
			15'h00002B94 : data <= 8'b00000000 ;
			15'h00002B95 : data <= 8'b00000000 ;
			15'h00002B96 : data <= 8'b00000000 ;
			15'h00002B97 : data <= 8'b00000000 ;
			15'h00002B98 : data <= 8'b00000000 ;
			15'h00002B99 : data <= 8'b00000000 ;
			15'h00002B9A : data <= 8'b00000000 ;
			15'h00002B9B : data <= 8'b00000000 ;
			15'h00002B9C : data <= 8'b00000000 ;
			15'h00002B9D : data <= 8'b00000000 ;
			15'h00002B9E : data <= 8'b00000000 ;
			15'h00002B9F : data <= 8'b00000000 ;
			15'h00002BA0 : data <= 8'b00000000 ;
			15'h00002BA1 : data <= 8'b00000000 ;
			15'h00002BA2 : data <= 8'b00000000 ;
			15'h00002BA3 : data <= 8'b00000000 ;
			15'h00002BA4 : data <= 8'b00000000 ;
			15'h00002BA5 : data <= 8'b00000000 ;
			15'h00002BA6 : data <= 8'b00000000 ;
			15'h00002BA7 : data <= 8'b00000000 ;
			15'h00002BA8 : data <= 8'b00000000 ;
			15'h00002BA9 : data <= 8'b00000000 ;
			15'h00002BAA : data <= 8'b00000000 ;
			15'h00002BAB : data <= 8'b00000000 ;
			15'h00002BAC : data <= 8'b00000000 ;
			15'h00002BAD : data <= 8'b00000000 ;
			15'h00002BAE : data <= 8'b00000000 ;
			15'h00002BAF : data <= 8'b00000000 ;
			15'h00002BB0 : data <= 8'b00000000 ;
			15'h00002BB1 : data <= 8'b00000000 ;
			15'h00002BB2 : data <= 8'b00000000 ;
			15'h00002BB3 : data <= 8'b00000000 ;
			15'h00002BB4 : data <= 8'b00000000 ;
			15'h00002BB5 : data <= 8'b00000000 ;
			15'h00002BB6 : data <= 8'b00000000 ;
			15'h00002BB7 : data <= 8'b00000000 ;
			15'h00002BB8 : data <= 8'b00000000 ;
			15'h00002BB9 : data <= 8'b00000000 ;
			15'h00002BBA : data <= 8'b00000000 ;
			15'h00002BBB : data <= 8'b00000000 ;
			15'h00002BBC : data <= 8'b00000000 ;
			15'h00002BBD : data <= 8'b00000000 ;
			15'h00002BBE : data <= 8'b00000000 ;
			15'h00002BBF : data <= 8'b00000000 ;
			15'h00002BC0 : data <= 8'b00000000 ;
			15'h00002BC1 : data <= 8'b00000000 ;
			15'h00002BC2 : data <= 8'b00000000 ;
			15'h00002BC3 : data <= 8'b00000000 ;
			15'h00002BC4 : data <= 8'b00000000 ;
			15'h00002BC5 : data <= 8'b00000000 ;
			15'h00002BC6 : data <= 8'b00000000 ;
			15'h00002BC7 : data <= 8'b00000000 ;
			15'h00002BC8 : data <= 8'b00000000 ;
			15'h00002BC9 : data <= 8'b00000000 ;
			15'h00002BCA : data <= 8'b00000000 ;
			15'h00002BCB : data <= 8'b00000000 ;
			15'h00002BCC : data <= 8'b00000000 ;
			15'h00002BCD : data <= 8'b00000000 ;
			15'h00002BCE : data <= 8'b00000000 ;
			15'h00002BCF : data <= 8'b00000000 ;
			15'h00002BD0 : data <= 8'b00000000 ;
			15'h00002BD1 : data <= 8'b00000000 ;
			15'h00002BD2 : data <= 8'b00000000 ;
			15'h00002BD3 : data <= 8'b00000000 ;
			15'h00002BD4 : data <= 8'b00000000 ;
			15'h00002BD5 : data <= 8'b00000000 ;
			15'h00002BD6 : data <= 8'b00000000 ;
			15'h00002BD7 : data <= 8'b00000000 ;
			15'h00002BD8 : data <= 8'b00000000 ;
			15'h00002BD9 : data <= 8'b00000000 ;
			15'h00002BDA : data <= 8'b00000000 ;
			15'h00002BDB : data <= 8'b00000000 ;
			15'h00002BDC : data <= 8'b00000000 ;
			15'h00002BDD : data <= 8'b00000000 ;
			15'h00002BDE : data <= 8'b00000000 ;
			15'h00002BDF : data <= 8'b00000000 ;
			15'h00002BE0 : data <= 8'b00000000 ;
			15'h00002BE1 : data <= 8'b00000000 ;
			15'h00002BE2 : data <= 8'b00000000 ;
			15'h00002BE3 : data <= 8'b00000000 ;
			15'h00002BE4 : data <= 8'b00000000 ;
			15'h00002BE5 : data <= 8'b00000000 ;
			15'h00002BE6 : data <= 8'b00000000 ;
			15'h00002BE7 : data <= 8'b00000000 ;
			15'h00002BE8 : data <= 8'b00000000 ;
			15'h00002BE9 : data <= 8'b00000000 ;
			15'h00002BEA : data <= 8'b00000000 ;
			15'h00002BEB : data <= 8'b00000000 ;
			15'h00002BEC : data <= 8'b00000000 ;
			15'h00002BED : data <= 8'b00000000 ;
			15'h00002BEE : data <= 8'b00000000 ;
			15'h00002BEF : data <= 8'b00000000 ;
			15'h00002BF0 : data <= 8'b00000000 ;
			15'h00002BF1 : data <= 8'b00000000 ;
			15'h00002BF2 : data <= 8'b00000000 ;
			15'h00002BF3 : data <= 8'b00000000 ;
			15'h00002BF4 : data <= 8'b00000000 ;
			15'h00002BF5 : data <= 8'b00000000 ;
			15'h00002BF6 : data <= 8'b00000000 ;
			15'h00002BF7 : data <= 8'b00000000 ;
			15'h00002BF8 : data <= 8'b00000000 ;
			15'h00002BF9 : data <= 8'b00000000 ;
			15'h00002BFA : data <= 8'b00000000 ;
			15'h00002BFB : data <= 8'b00000000 ;
			15'h00002BFC : data <= 8'b00000000 ;
			15'h00002BFD : data <= 8'b00000000 ;
			15'h00002BFE : data <= 8'b00000000 ;
			15'h00002BFF : data <= 8'b00000000 ;
			15'h00002C00 : data <= 8'b00000000 ;
			15'h00002C01 : data <= 8'b00000000 ;
			15'h00002C02 : data <= 8'b00000000 ;
			15'h00002C03 : data <= 8'b00000000 ;
			15'h00002C04 : data <= 8'b00000000 ;
			15'h00002C05 : data <= 8'b00000000 ;
			15'h00002C06 : data <= 8'b00000000 ;
			15'h00002C07 : data <= 8'b00000000 ;
			15'h00002C08 : data <= 8'b00000000 ;
			15'h00002C09 : data <= 8'b00000000 ;
			15'h00002C0A : data <= 8'b00000000 ;
			15'h00002C0B : data <= 8'b00000000 ;
			15'h00002C0C : data <= 8'b00000000 ;
			15'h00002C0D : data <= 8'b00000000 ;
			15'h00002C0E : data <= 8'b00000000 ;
			15'h00002C0F : data <= 8'b00000000 ;
			15'h00002C10 : data <= 8'b00000000 ;
			15'h00002C11 : data <= 8'b00000000 ;
			15'h00002C12 : data <= 8'b00000000 ;
			15'h00002C13 : data <= 8'b00000000 ;
			15'h00002C14 : data <= 8'b00000000 ;
			15'h00002C15 : data <= 8'b00000000 ;
			15'h00002C16 : data <= 8'b00000000 ;
			15'h00002C17 : data <= 8'b00000000 ;
			15'h00002C18 : data <= 8'b00000000 ;
			15'h00002C19 : data <= 8'b00000000 ;
			15'h00002C1A : data <= 8'b00000000 ;
			15'h00002C1B : data <= 8'b00000000 ;
			15'h00002C1C : data <= 8'b00000000 ;
			15'h00002C1D : data <= 8'b00000000 ;
			15'h00002C1E : data <= 8'b00000000 ;
			15'h00002C1F : data <= 8'b00000000 ;
			15'h00002C20 : data <= 8'b00000000 ;
			15'h00002C21 : data <= 8'b00000000 ;
			15'h00002C22 : data <= 8'b00000000 ;
			15'h00002C23 : data <= 8'b00000000 ;
			15'h00002C24 : data <= 8'b00000000 ;
			15'h00002C25 : data <= 8'b00000000 ;
			15'h00002C26 : data <= 8'b00000000 ;
			15'h00002C27 : data <= 8'b00000000 ;
			15'h00002C28 : data <= 8'b00000000 ;
			15'h00002C29 : data <= 8'b00000000 ;
			15'h00002C2A : data <= 8'b00000000 ;
			15'h00002C2B : data <= 8'b00000000 ;
			15'h00002C2C : data <= 8'b00000000 ;
			15'h00002C2D : data <= 8'b00000000 ;
			15'h00002C2E : data <= 8'b00000000 ;
			15'h00002C2F : data <= 8'b00000000 ;
			15'h00002C30 : data <= 8'b00000000 ;
			15'h00002C31 : data <= 8'b00000000 ;
			15'h00002C32 : data <= 8'b00000000 ;
			15'h00002C33 : data <= 8'b00000000 ;
			15'h00002C34 : data <= 8'b00000000 ;
			15'h00002C35 : data <= 8'b00000000 ;
			15'h00002C36 : data <= 8'b00000000 ;
			15'h00002C37 : data <= 8'b00000000 ;
			15'h00002C38 : data <= 8'b00000000 ;
			15'h00002C39 : data <= 8'b00000000 ;
			15'h00002C3A : data <= 8'b00000000 ;
			15'h00002C3B : data <= 8'b00000000 ;
			15'h00002C3C : data <= 8'b00000000 ;
			15'h00002C3D : data <= 8'b00000000 ;
			15'h00002C3E : data <= 8'b00000000 ;
			15'h00002C3F : data <= 8'b00000000 ;
			15'h00002C40 : data <= 8'b00000000 ;
			15'h00002C41 : data <= 8'b00000000 ;
			15'h00002C42 : data <= 8'b00000000 ;
			15'h00002C43 : data <= 8'b00000000 ;
			15'h00002C44 : data <= 8'b00000000 ;
			15'h00002C45 : data <= 8'b00000000 ;
			15'h00002C46 : data <= 8'b00000000 ;
			15'h00002C47 : data <= 8'b00000000 ;
			15'h00002C48 : data <= 8'b00000000 ;
			15'h00002C49 : data <= 8'b00000000 ;
			15'h00002C4A : data <= 8'b00000000 ;
			15'h00002C4B : data <= 8'b00000000 ;
			15'h00002C4C : data <= 8'b00000000 ;
			15'h00002C4D : data <= 8'b00000000 ;
			15'h00002C4E : data <= 8'b00000000 ;
			15'h00002C4F : data <= 8'b00000000 ;
			15'h00002C50 : data <= 8'b00000000 ;
			15'h00002C51 : data <= 8'b00000000 ;
			15'h00002C52 : data <= 8'b00000000 ;
			15'h00002C53 : data <= 8'b00000000 ;
			15'h00002C54 : data <= 8'b00000000 ;
			15'h00002C55 : data <= 8'b00000000 ;
			15'h00002C56 : data <= 8'b00000000 ;
			15'h00002C57 : data <= 8'b00000000 ;
			15'h00002C58 : data <= 8'b00000000 ;
			15'h00002C59 : data <= 8'b00000000 ;
			15'h00002C5A : data <= 8'b00000000 ;
			15'h00002C5B : data <= 8'b00000000 ;
			15'h00002C5C : data <= 8'b00000000 ;
			15'h00002C5D : data <= 8'b00000000 ;
			15'h00002C5E : data <= 8'b00000000 ;
			15'h00002C5F : data <= 8'b00000000 ;
			15'h00002C60 : data <= 8'b00000000 ;
			15'h00002C61 : data <= 8'b00000000 ;
			15'h00002C62 : data <= 8'b00000000 ;
			15'h00002C63 : data <= 8'b00000000 ;
			15'h00002C64 : data <= 8'b00000000 ;
			15'h00002C65 : data <= 8'b00000000 ;
			15'h00002C66 : data <= 8'b00000000 ;
			15'h00002C67 : data <= 8'b00000000 ;
			15'h00002C68 : data <= 8'b00000000 ;
			15'h00002C69 : data <= 8'b00000000 ;
			15'h00002C6A : data <= 8'b00000000 ;
			15'h00002C6B : data <= 8'b00000000 ;
			15'h00002C6C : data <= 8'b00000000 ;
			15'h00002C6D : data <= 8'b00000000 ;
			15'h00002C6E : data <= 8'b00000000 ;
			15'h00002C6F : data <= 8'b00000000 ;
			15'h00002C70 : data <= 8'b00000000 ;
			15'h00002C71 : data <= 8'b00000000 ;
			15'h00002C72 : data <= 8'b00000000 ;
			15'h00002C73 : data <= 8'b00000000 ;
			15'h00002C74 : data <= 8'b00000000 ;
			15'h00002C75 : data <= 8'b00000000 ;
			15'h00002C76 : data <= 8'b00000000 ;
			15'h00002C77 : data <= 8'b00000000 ;
			15'h00002C78 : data <= 8'b00000000 ;
			15'h00002C79 : data <= 8'b00000000 ;
			15'h00002C7A : data <= 8'b00000000 ;
			15'h00002C7B : data <= 8'b00000000 ;
			15'h00002C7C : data <= 8'b00000000 ;
			15'h00002C7D : data <= 8'b00000000 ;
			15'h00002C7E : data <= 8'b00000000 ;
			15'h00002C7F : data <= 8'b00000000 ;
			15'h00002C80 : data <= 8'b00000000 ;
			15'h00002C81 : data <= 8'b00000000 ;
			15'h00002C82 : data <= 8'b00000000 ;
			15'h00002C83 : data <= 8'b00000000 ;
			15'h00002C84 : data <= 8'b00000000 ;
			15'h00002C85 : data <= 8'b00000000 ;
			15'h00002C86 : data <= 8'b00000000 ;
			15'h00002C87 : data <= 8'b00000000 ;
			15'h00002C88 : data <= 8'b00000000 ;
			15'h00002C89 : data <= 8'b00000000 ;
			15'h00002C8A : data <= 8'b00000000 ;
			15'h00002C8B : data <= 8'b00000000 ;
			15'h00002C8C : data <= 8'b00000000 ;
			15'h00002C8D : data <= 8'b00000000 ;
			15'h00002C8E : data <= 8'b00000000 ;
			15'h00002C8F : data <= 8'b00000000 ;
			15'h00002C90 : data <= 8'b00000000 ;
			15'h00002C91 : data <= 8'b00000000 ;
			15'h00002C92 : data <= 8'b00000000 ;
			15'h00002C93 : data <= 8'b00000000 ;
			15'h00002C94 : data <= 8'b00000000 ;
			15'h00002C95 : data <= 8'b00000000 ;
			15'h00002C96 : data <= 8'b00000000 ;
			15'h00002C97 : data <= 8'b00000000 ;
			15'h00002C98 : data <= 8'b00000000 ;
			15'h00002C99 : data <= 8'b00000000 ;
			15'h00002C9A : data <= 8'b00000000 ;
			15'h00002C9B : data <= 8'b00000000 ;
			15'h00002C9C : data <= 8'b00000000 ;
			15'h00002C9D : data <= 8'b00000000 ;
			15'h00002C9E : data <= 8'b00000000 ;
			15'h00002C9F : data <= 8'b00000000 ;
			15'h00002CA0 : data <= 8'b00000000 ;
			15'h00002CA1 : data <= 8'b00000000 ;
			15'h00002CA2 : data <= 8'b00000000 ;
			15'h00002CA3 : data <= 8'b00000000 ;
			15'h00002CA4 : data <= 8'b00000000 ;
			15'h00002CA5 : data <= 8'b00000000 ;
			15'h00002CA6 : data <= 8'b00000000 ;
			15'h00002CA7 : data <= 8'b00000000 ;
			15'h00002CA8 : data <= 8'b00000000 ;
			15'h00002CA9 : data <= 8'b00000000 ;
			15'h00002CAA : data <= 8'b00000000 ;
			15'h00002CAB : data <= 8'b00000000 ;
			15'h00002CAC : data <= 8'b00000000 ;
			15'h00002CAD : data <= 8'b00000000 ;
			15'h00002CAE : data <= 8'b00000000 ;
			15'h00002CAF : data <= 8'b00000000 ;
			15'h00002CB0 : data <= 8'b00000000 ;
			15'h00002CB1 : data <= 8'b00000000 ;
			15'h00002CB2 : data <= 8'b00000000 ;
			15'h00002CB3 : data <= 8'b00000000 ;
			15'h00002CB4 : data <= 8'b00000000 ;
			15'h00002CB5 : data <= 8'b00000000 ;
			15'h00002CB6 : data <= 8'b00000000 ;
			15'h00002CB7 : data <= 8'b00000000 ;
			15'h00002CB8 : data <= 8'b00000000 ;
			15'h00002CB9 : data <= 8'b00000000 ;
			15'h00002CBA : data <= 8'b00000000 ;
			15'h00002CBB : data <= 8'b00000000 ;
			15'h00002CBC : data <= 8'b00000000 ;
			15'h00002CBD : data <= 8'b00000000 ;
			15'h00002CBE : data <= 8'b00000000 ;
			15'h00002CBF : data <= 8'b00000000 ;
			15'h00002CC0 : data <= 8'b00000000 ;
			15'h00002CC1 : data <= 8'b00000000 ;
			15'h00002CC2 : data <= 8'b00000000 ;
			15'h00002CC3 : data <= 8'b00000000 ;
			15'h00002CC4 : data <= 8'b00000000 ;
			15'h00002CC5 : data <= 8'b00000000 ;
			15'h00002CC6 : data <= 8'b00000000 ;
			15'h00002CC7 : data <= 8'b00000000 ;
			15'h00002CC8 : data <= 8'b00000000 ;
			15'h00002CC9 : data <= 8'b00000000 ;
			15'h00002CCA : data <= 8'b00000000 ;
			15'h00002CCB : data <= 8'b00000000 ;
			15'h00002CCC : data <= 8'b00000000 ;
			15'h00002CCD : data <= 8'b00000000 ;
			15'h00002CCE : data <= 8'b00000000 ;
			15'h00002CCF : data <= 8'b00000000 ;
			15'h00002CD0 : data <= 8'b00000000 ;
			15'h00002CD1 : data <= 8'b00000000 ;
			15'h00002CD2 : data <= 8'b00000000 ;
			15'h00002CD3 : data <= 8'b00000000 ;
			15'h00002CD4 : data <= 8'b00000000 ;
			15'h00002CD5 : data <= 8'b00000000 ;
			15'h00002CD6 : data <= 8'b00000000 ;
			15'h00002CD7 : data <= 8'b00000000 ;
			15'h00002CD8 : data <= 8'b00000000 ;
			15'h00002CD9 : data <= 8'b00000000 ;
			15'h00002CDA : data <= 8'b00000000 ;
			15'h00002CDB : data <= 8'b00000000 ;
			15'h00002CDC : data <= 8'b00000000 ;
			15'h00002CDD : data <= 8'b00000000 ;
			15'h00002CDE : data <= 8'b00000000 ;
			15'h00002CDF : data <= 8'b00000000 ;
			15'h00002CE0 : data <= 8'b00000000 ;
			15'h00002CE1 : data <= 8'b00000000 ;
			15'h00002CE2 : data <= 8'b00000000 ;
			15'h00002CE3 : data <= 8'b00000000 ;
			15'h00002CE4 : data <= 8'b00000000 ;
			15'h00002CE5 : data <= 8'b00000000 ;
			15'h00002CE6 : data <= 8'b00000000 ;
			15'h00002CE7 : data <= 8'b00000000 ;
			15'h00002CE8 : data <= 8'b00000000 ;
			15'h00002CE9 : data <= 8'b00000000 ;
			15'h00002CEA : data <= 8'b00000000 ;
			15'h00002CEB : data <= 8'b00000000 ;
			15'h00002CEC : data <= 8'b00000000 ;
			15'h00002CED : data <= 8'b00000000 ;
			15'h00002CEE : data <= 8'b00000000 ;
			15'h00002CEF : data <= 8'b00000000 ;
			15'h00002CF0 : data <= 8'b00000000 ;
			15'h00002CF1 : data <= 8'b00000000 ;
			15'h00002CF2 : data <= 8'b00000000 ;
			15'h00002CF3 : data <= 8'b00000000 ;
			15'h00002CF4 : data <= 8'b00000000 ;
			15'h00002CF5 : data <= 8'b00000000 ;
			15'h00002CF6 : data <= 8'b00000000 ;
			15'h00002CF7 : data <= 8'b00000000 ;
			15'h00002CF8 : data <= 8'b00000000 ;
			15'h00002CF9 : data <= 8'b00000000 ;
			15'h00002CFA : data <= 8'b00000000 ;
			15'h00002CFB : data <= 8'b00000000 ;
			15'h00002CFC : data <= 8'b00000000 ;
			15'h00002CFD : data <= 8'b00000000 ;
			15'h00002CFE : data <= 8'b00000000 ;
			15'h00002CFF : data <= 8'b00000000 ;
			15'h00002D00 : data <= 8'b00000000 ;
			15'h00002D01 : data <= 8'b00000000 ;
			15'h00002D02 : data <= 8'b00000000 ;
			15'h00002D03 : data <= 8'b00000000 ;
			15'h00002D04 : data <= 8'b00000000 ;
			15'h00002D05 : data <= 8'b00000000 ;
			15'h00002D06 : data <= 8'b00000000 ;
			15'h00002D07 : data <= 8'b00000000 ;
			15'h00002D08 : data <= 8'b00000000 ;
			15'h00002D09 : data <= 8'b00000000 ;
			15'h00002D0A : data <= 8'b00000000 ;
			15'h00002D0B : data <= 8'b00000000 ;
			15'h00002D0C : data <= 8'b00000000 ;
			15'h00002D0D : data <= 8'b00000000 ;
			15'h00002D0E : data <= 8'b00000000 ;
			15'h00002D0F : data <= 8'b00000000 ;
			15'h00002D10 : data <= 8'b00000000 ;
			15'h00002D11 : data <= 8'b00000000 ;
			15'h00002D12 : data <= 8'b00000000 ;
			15'h00002D13 : data <= 8'b00000000 ;
			15'h00002D14 : data <= 8'b00000000 ;
			15'h00002D15 : data <= 8'b00000000 ;
			15'h00002D16 : data <= 8'b00000000 ;
			15'h00002D17 : data <= 8'b00000000 ;
			15'h00002D18 : data <= 8'b00000000 ;
			15'h00002D19 : data <= 8'b00000000 ;
			15'h00002D1A : data <= 8'b00000000 ;
			15'h00002D1B : data <= 8'b00000000 ;
			15'h00002D1C : data <= 8'b00000000 ;
			15'h00002D1D : data <= 8'b00000000 ;
			15'h00002D1E : data <= 8'b00000000 ;
			15'h00002D1F : data <= 8'b00000000 ;
			15'h00002D20 : data <= 8'b00000000 ;
			15'h00002D21 : data <= 8'b00000000 ;
			15'h00002D22 : data <= 8'b00000000 ;
			15'h00002D23 : data <= 8'b00000000 ;
			15'h00002D24 : data <= 8'b00000000 ;
			15'h00002D25 : data <= 8'b00000000 ;
			15'h00002D26 : data <= 8'b00000000 ;
			15'h00002D27 : data <= 8'b00000000 ;
			15'h00002D28 : data <= 8'b00000000 ;
			15'h00002D29 : data <= 8'b00000000 ;
			15'h00002D2A : data <= 8'b00000000 ;
			15'h00002D2B : data <= 8'b00000000 ;
			15'h00002D2C : data <= 8'b00000000 ;
			15'h00002D2D : data <= 8'b00000000 ;
			15'h00002D2E : data <= 8'b00000000 ;
			15'h00002D2F : data <= 8'b00000000 ;
			15'h00002D30 : data <= 8'b00000000 ;
			15'h00002D31 : data <= 8'b00000000 ;
			15'h00002D32 : data <= 8'b00000000 ;
			15'h00002D33 : data <= 8'b00000000 ;
			15'h00002D34 : data <= 8'b00000000 ;
			15'h00002D35 : data <= 8'b00000000 ;
			15'h00002D36 : data <= 8'b00000000 ;
			15'h00002D37 : data <= 8'b00000000 ;
			15'h00002D38 : data <= 8'b00000000 ;
			15'h00002D39 : data <= 8'b00000000 ;
			15'h00002D3A : data <= 8'b00000000 ;
			15'h00002D3B : data <= 8'b00000000 ;
			15'h00002D3C : data <= 8'b00000000 ;
			15'h00002D3D : data <= 8'b00000000 ;
			15'h00002D3E : data <= 8'b00000000 ;
			15'h00002D3F : data <= 8'b00000000 ;
			15'h00002D40 : data <= 8'b00000000 ;
			15'h00002D41 : data <= 8'b00000000 ;
			15'h00002D42 : data <= 8'b00000000 ;
			15'h00002D43 : data <= 8'b00000000 ;
			15'h00002D44 : data <= 8'b00000000 ;
			15'h00002D45 : data <= 8'b00000000 ;
			15'h00002D46 : data <= 8'b00000000 ;
			15'h00002D47 : data <= 8'b00000000 ;
			15'h00002D48 : data <= 8'b00000000 ;
			15'h00002D49 : data <= 8'b00000000 ;
			15'h00002D4A : data <= 8'b00000000 ;
			15'h00002D4B : data <= 8'b00000000 ;
			15'h00002D4C : data <= 8'b00000000 ;
			15'h00002D4D : data <= 8'b00000000 ;
			15'h00002D4E : data <= 8'b00000000 ;
			15'h00002D4F : data <= 8'b00000000 ;
			15'h00002D50 : data <= 8'b00000000 ;
			15'h00002D51 : data <= 8'b00000000 ;
			15'h00002D52 : data <= 8'b00000000 ;
			15'h00002D53 : data <= 8'b00000000 ;
			15'h00002D54 : data <= 8'b00000000 ;
			15'h00002D55 : data <= 8'b00000000 ;
			15'h00002D56 : data <= 8'b00000000 ;
			15'h00002D57 : data <= 8'b00000000 ;
			15'h00002D58 : data <= 8'b00000000 ;
			15'h00002D59 : data <= 8'b00000000 ;
			15'h00002D5A : data <= 8'b00000000 ;
			15'h00002D5B : data <= 8'b00000000 ;
			15'h00002D5C : data <= 8'b00000000 ;
			15'h00002D5D : data <= 8'b00000000 ;
			15'h00002D5E : data <= 8'b00000000 ;
			15'h00002D5F : data <= 8'b00000000 ;
			15'h00002D60 : data <= 8'b00000000 ;
			15'h00002D61 : data <= 8'b00000000 ;
			15'h00002D62 : data <= 8'b00000000 ;
			15'h00002D63 : data <= 8'b00000000 ;
			15'h00002D64 : data <= 8'b00000000 ;
			15'h00002D65 : data <= 8'b00000000 ;
			15'h00002D66 : data <= 8'b00000000 ;
			15'h00002D67 : data <= 8'b00000000 ;
			15'h00002D68 : data <= 8'b00000000 ;
			15'h00002D69 : data <= 8'b00000000 ;
			15'h00002D6A : data <= 8'b00000000 ;
			15'h00002D6B : data <= 8'b00000000 ;
			15'h00002D6C : data <= 8'b00000000 ;
			15'h00002D6D : data <= 8'b00000000 ;
			15'h00002D6E : data <= 8'b00000000 ;
			15'h00002D6F : data <= 8'b00000000 ;
			15'h00002D70 : data <= 8'b00000000 ;
			15'h00002D71 : data <= 8'b00000000 ;
			15'h00002D72 : data <= 8'b00000000 ;
			15'h00002D73 : data <= 8'b00000000 ;
			15'h00002D74 : data <= 8'b00000000 ;
			15'h00002D75 : data <= 8'b00000000 ;
			15'h00002D76 : data <= 8'b00000000 ;
			15'h00002D77 : data <= 8'b00000000 ;
			15'h00002D78 : data <= 8'b00000000 ;
			15'h00002D79 : data <= 8'b00000000 ;
			15'h00002D7A : data <= 8'b00000000 ;
			15'h00002D7B : data <= 8'b00000000 ;
			15'h00002D7C : data <= 8'b00000000 ;
			15'h00002D7D : data <= 8'b00000000 ;
			15'h00002D7E : data <= 8'b00000000 ;
			15'h00002D7F : data <= 8'b00000000 ;
			15'h00002D80 : data <= 8'b00000000 ;
			15'h00002D81 : data <= 8'b00000000 ;
			15'h00002D82 : data <= 8'b00000000 ;
			15'h00002D83 : data <= 8'b00000000 ;
			15'h00002D84 : data <= 8'b00000000 ;
			15'h00002D85 : data <= 8'b00000000 ;
			15'h00002D86 : data <= 8'b00000000 ;
			15'h00002D87 : data <= 8'b00000000 ;
			15'h00002D88 : data <= 8'b00000000 ;
			15'h00002D89 : data <= 8'b00000000 ;
			15'h00002D8A : data <= 8'b00000000 ;
			15'h00002D8B : data <= 8'b00000000 ;
			15'h00002D8C : data <= 8'b00000000 ;
			15'h00002D8D : data <= 8'b00000000 ;
			15'h00002D8E : data <= 8'b00000000 ;
			15'h00002D8F : data <= 8'b00000000 ;
			15'h00002D90 : data <= 8'b00000000 ;
			15'h00002D91 : data <= 8'b00000000 ;
			15'h00002D92 : data <= 8'b00000000 ;
			15'h00002D93 : data <= 8'b00000000 ;
			15'h00002D94 : data <= 8'b00000000 ;
			15'h00002D95 : data <= 8'b00000000 ;
			15'h00002D96 : data <= 8'b00000000 ;
			15'h00002D97 : data <= 8'b00000000 ;
			15'h00002D98 : data <= 8'b00000000 ;
			15'h00002D99 : data <= 8'b00000000 ;
			15'h00002D9A : data <= 8'b00000000 ;
			15'h00002D9B : data <= 8'b00000000 ;
			15'h00002D9C : data <= 8'b00000000 ;
			15'h00002D9D : data <= 8'b00000000 ;
			15'h00002D9E : data <= 8'b00000000 ;
			15'h00002D9F : data <= 8'b00000000 ;
			15'h00002DA0 : data <= 8'b00000000 ;
			15'h00002DA1 : data <= 8'b00000000 ;
			15'h00002DA2 : data <= 8'b00000000 ;
			15'h00002DA3 : data <= 8'b00000000 ;
			15'h00002DA4 : data <= 8'b00000000 ;
			15'h00002DA5 : data <= 8'b00000000 ;
			15'h00002DA6 : data <= 8'b00000000 ;
			15'h00002DA7 : data <= 8'b00000000 ;
			15'h00002DA8 : data <= 8'b00000000 ;
			15'h00002DA9 : data <= 8'b00000000 ;
			15'h00002DAA : data <= 8'b00000000 ;
			15'h00002DAB : data <= 8'b00000000 ;
			15'h00002DAC : data <= 8'b00000000 ;
			15'h00002DAD : data <= 8'b00000000 ;
			15'h00002DAE : data <= 8'b00000000 ;
			15'h00002DAF : data <= 8'b00000000 ;
			15'h00002DB0 : data <= 8'b00000000 ;
			15'h00002DB1 : data <= 8'b00000000 ;
			15'h00002DB2 : data <= 8'b00000000 ;
			15'h00002DB3 : data <= 8'b00000000 ;
			15'h00002DB4 : data <= 8'b00000000 ;
			15'h00002DB5 : data <= 8'b00000000 ;
			15'h00002DB6 : data <= 8'b00000000 ;
			15'h00002DB7 : data <= 8'b00000000 ;
			15'h00002DB8 : data <= 8'b00000000 ;
			15'h00002DB9 : data <= 8'b00000000 ;
			15'h00002DBA : data <= 8'b00000000 ;
			15'h00002DBB : data <= 8'b00000000 ;
			15'h00002DBC : data <= 8'b00000000 ;
			15'h00002DBD : data <= 8'b00000000 ;
			15'h00002DBE : data <= 8'b00000000 ;
			15'h00002DBF : data <= 8'b00000000 ;
			15'h00002DC0 : data <= 8'b00000000 ;
			15'h00002DC1 : data <= 8'b00000000 ;
			15'h00002DC2 : data <= 8'b00000000 ;
			15'h00002DC3 : data <= 8'b00000000 ;
			15'h00002DC4 : data <= 8'b00000000 ;
			15'h00002DC5 : data <= 8'b00000000 ;
			15'h00002DC6 : data <= 8'b00000000 ;
			15'h00002DC7 : data <= 8'b00000000 ;
			15'h00002DC8 : data <= 8'b00000000 ;
			15'h00002DC9 : data <= 8'b00000000 ;
			15'h00002DCA : data <= 8'b00000000 ;
			15'h00002DCB : data <= 8'b00000000 ;
			15'h00002DCC : data <= 8'b00000000 ;
			15'h00002DCD : data <= 8'b00000000 ;
			15'h00002DCE : data <= 8'b00000000 ;
			15'h00002DCF : data <= 8'b00000000 ;
			15'h00002DD0 : data <= 8'b00000000 ;
			15'h00002DD1 : data <= 8'b00000000 ;
			15'h00002DD2 : data <= 8'b00000000 ;
			15'h00002DD3 : data <= 8'b00000000 ;
			15'h00002DD4 : data <= 8'b00000000 ;
			15'h00002DD5 : data <= 8'b00000000 ;
			15'h00002DD6 : data <= 8'b00000000 ;
			15'h00002DD7 : data <= 8'b00000000 ;
			15'h00002DD8 : data <= 8'b00000000 ;
			15'h00002DD9 : data <= 8'b00000000 ;
			15'h00002DDA : data <= 8'b00000000 ;
			15'h00002DDB : data <= 8'b00000000 ;
			15'h00002DDC : data <= 8'b00000000 ;
			15'h00002DDD : data <= 8'b00000000 ;
			15'h00002DDE : data <= 8'b00000000 ;
			15'h00002DDF : data <= 8'b00000000 ;
			15'h00002DE0 : data <= 8'b00000000 ;
			15'h00002DE1 : data <= 8'b00000000 ;
			15'h00002DE2 : data <= 8'b00000000 ;
			15'h00002DE3 : data <= 8'b00000000 ;
			15'h00002DE4 : data <= 8'b00000000 ;
			15'h00002DE5 : data <= 8'b00000000 ;
			15'h00002DE6 : data <= 8'b00000000 ;
			15'h00002DE7 : data <= 8'b00000000 ;
			15'h00002DE8 : data <= 8'b00000000 ;
			15'h00002DE9 : data <= 8'b00000000 ;
			15'h00002DEA : data <= 8'b00000000 ;
			15'h00002DEB : data <= 8'b00000000 ;
			15'h00002DEC : data <= 8'b00000000 ;
			15'h00002DED : data <= 8'b00000000 ;
			15'h00002DEE : data <= 8'b00000000 ;
			15'h00002DEF : data <= 8'b00000000 ;
			15'h00002DF0 : data <= 8'b00000000 ;
			15'h00002DF1 : data <= 8'b00000000 ;
			15'h00002DF2 : data <= 8'b00000000 ;
			15'h00002DF3 : data <= 8'b00000000 ;
			15'h00002DF4 : data <= 8'b00000000 ;
			15'h00002DF5 : data <= 8'b00000000 ;
			15'h00002DF6 : data <= 8'b00000000 ;
			15'h00002DF7 : data <= 8'b00000000 ;
			15'h00002DF8 : data <= 8'b00000000 ;
			15'h00002DF9 : data <= 8'b00000000 ;
			15'h00002DFA : data <= 8'b00000000 ;
			15'h00002DFB : data <= 8'b00000000 ;
			15'h00002DFC : data <= 8'b00000000 ;
			15'h00002DFD : data <= 8'b00000000 ;
			15'h00002DFE : data <= 8'b00000000 ;
			15'h00002DFF : data <= 8'b00000000 ;
			15'h00002E00 : data <= 8'b00000000 ;
			15'h00002E01 : data <= 8'b00000000 ;
			15'h00002E02 : data <= 8'b00000000 ;
			15'h00002E03 : data <= 8'b00000000 ;
			15'h00002E04 : data <= 8'b00000000 ;
			15'h00002E05 : data <= 8'b00000000 ;
			15'h00002E06 : data <= 8'b00000000 ;
			15'h00002E07 : data <= 8'b00000000 ;
			15'h00002E08 : data <= 8'b00000000 ;
			15'h00002E09 : data <= 8'b00000000 ;
			15'h00002E0A : data <= 8'b00000000 ;
			15'h00002E0B : data <= 8'b00000000 ;
			15'h00002E0C : data <= 8'b00000000 ;
			15'h00002E0D : data <= 8'b00000000 ;
			15'h00002E0E : data <= 8'b00000000 ;
			15'h00002E0F : data <= 8'b00000000 ;
			15'h00002E10 : data <= 8'b00000000 ;
			15'h00002E11 : data <= 8'b00000000 ;
			15'h00002E12 : data <= 8'b00000000 ;
			15'h00002E13 : data <= 8'b00000000 ;
			15'h00002E14 : data <= 8'b00000000 ;
			15'h00002E15 : data <= 8'b00000000 ;
			15'h00002E16 : data <= 8'b00000000 ;
			15'h00002E17 : data <= 8'b00000000 ;
			15'h00002E18 : data <= 8'b00000000 ;
			15'h00002E19 : data <= 8'b00000000 ;
			15'h00002E1A : data <= 8'b00000000 ;
			15'h00002E1B : data <= 8'b00000000 ;
			15'h00002E1C : data <= 8'b00000000 ;
			15'h00002E1D : data <= 8'b00000000 ;
			15'h00002E1E : data <= 8'b00000000 ;
			15'h00002E1F : data <= 8'b00000000 ;
			15'h00002E20 : data <= 8'b00000000 ;
			15'h00002E21 : data <= 8'b00000000 ;
			15'h00002E22 : data <= 8'b00000000 ;
			15'h00002E23 : data <= 8'b00000000 ;
			15'h00002E24 : data <= 8'b00000000 ;
			15'h00002E25 : data <= 8'b00000000 ;
			15'h00002E26 : data <= 8'b00000000 ;
			15'h00002E27 : data <= 8'b00000000 ;
			15'h00002E28 : data <= 8'b00000000 ;
			15'h00002E29 : data <= 8'b00000000 ;
			15'h00002E2A : data <= 8'b00000000 ;
			15'h00002E2B : data <= 8'b00000000 ;
			15'h00002E2C : data <= 8'b00000000 ;
			15'h00002E2D : data <= 8'b00000000 ;
			15'h00002E2E : data <= 8'b00000000 ;
			15'h00002E2F : data <= 8'b00000000 ;
			15'h00002E30 : data <= 8'b00000000 ;
			15'h00002E31 : data <= 8'b00000000 ;
			15'h00002E32 : data <= 8'b00000000 ;
			15'h00002E33 : data <= 8'b00000000 ;
			15'h00002E34 : data <= 8'b00000000 ;
			15'h00002E35 : data <= 8'b00000000 ;
			15'h00002E36 : data <= 8'b00000000 ;
			15'h00002E37 : data <= 8'b00000000 ;
			15'h00002E38 : data <= 8'b00000000 ;
			15'h00002E39 : data <= 8'b00000000 ;
			15'h00002E3A : data <= 8'b00000000 ;
			15'h00002E3B : data <= 8'b00000000 ;
			15'h00002E3C : data <= 8'b00000000 ;
			15'h00002E3D : data <= 8'b00000000 ;
			15'h00002E3E : data <= 8'b00000000 ;
			15'h00002E3F : data <= 8'b00000000 ;
			15'h00002E40 : data <= 8'b00000000 ;
			15'h00002E41 : data <= 8'b00000000 ;
			15'h00002E42 : data <= 8'b00000000 ;
			15'h00002E43 : data <= 8'b00000000 ;
			15'h00002E44 : data <= 8'b00000000 ;
			15'h00002E45 : data <= 8'b00000000 ;
			15'h00002E46 : data <= 8'b00000000 ;
			15'h00002E47 : data <= 8'b00000000 ;
			15'h00002E48 : data <= 8'b00000000 ;
			15'h00002E49 : data <= 8'b00000000 ;
			15'h00002E4A : data <= 8'b00000000 ;
			15'h00002E4B : data <= 8'b00000000 ;
			15'h00002E4C : data <= 8'b00000000 ;
			15'h00002E4D : data <= 8'b00000000 ;
			15'h00002E4E : data <= 8'b00000000 ;
			15'h00002E4F : data <= 8'b00000000 ;
			15'h00002E50 : data <= 8'b00000000 ;
			15'h00002E51 : data <= 8'b00000000 ;
			15'h00002E52 : data <= 8'b00000000 ;
			15'h00002E53 : data <= 8'b00000000 ;
			15'h00002E54 : data <= 8'b00000000 ;
			15'h00002E55 : data <= 8'b00000000 ;
			15'h00002E56 : data <= 8'b00000000 ;
			15'h00002E57 : data <= 8'b00000000 ;
			15'h00002E58 : data <= 8'b00000000 ;
			15'h00002E59 : data <= 8'b00000000 ;
			15'h00002E5A : data <= 8'b00000000 ;
			15'h00002E5B : data <= 8'b00000000 ;
			15'h00002E5C : data <= 8'b00000000 ;
			15'h00002E5D : data <= 8'b00000000 ;
			15'h00002E5E : data <= 8'b00000000 ;
			15'h00002E5F : data <= 8'b00000000 ;
			15'h00002E60 : data <= 8'b00000000 ;
			15'h00002E61 : data <= 8'b00000000 ;
			15'h00002E62 : data <= 8'b00000000 ;
			15'h00002E63 : data <= 8'b00000000 ;
			15'h00002E64 : data <= 8'b00000000 ;
			15'h00002E65 : data <= 8'b00000000 ;
			15'h00002E66 : data <= 8'b00000000 ;
			15'h00002E67 : data <= 8'b00000000 ;
			15'h00002E68 : data <= 8'b00000000 ;
			15'h00002E69 : data <= 8'b00000000 ;
			15'h00002E6A : data <= 8'b00000000 ;
			15'h00002E6B : data <= 8'b00000000 ;
			15'h00002E6C : data <= 8'b00000000 ;
			15'h00002E6D : data <= 8'b00000000 ;
			15'h00002E6E : data <= 8'b00000000 ;
			15'h00002E6F : data <= 8'b00000000 ;
			15'h00002E70 : data <= 8'b00000000 ;
			15'h00002E71 : data <= 8'b00000000 ;
			15'h00002E72 : data <= 8'b00000000 ;
			15'h00002E73 : data <= 8'b00000000 ;
			15'h00002E74 : data <= 8'b00000000 ;
			15'h00002E75 : data <= 8'b00000000 ;
			15'h00002E76 : data <= 8'b00000000 ;
			15'h00002E77 : data <= 8'b00000000 ;
			15'h00002E78 : data <= 8'b00000000 ;
			15'h00002E79 : data <= 8'b00000000 ;
			15'h00002E7A : data <= 8'b00000000 ;
			15'h00002E7B : data <= 8'b00000000 ;
			15'h00002E7C : data <= 8'b00000000 ;
			15'h00002E7D : data <= 8'b00000000 ;
			15'h00002E7E : data <= 8'b00000000 ;
			15'h00002E7F : data <= 8'b00000000 ;
			15'h00002E80 : data <= 8'b00000000 ;
			15'h00002E81 : data <= 8'b00000000 ;
			15'h00002E82 : data <= 8'b00000000 ;
			15'h00002E83 : data <= 8'b00000000 ;
			15'h00002E84 : data <= 8'b00000000 ;
			15'h00002E85 : data <= 8'b00000000 ;
			15'h00002E86 : data <= 8'b00000000 ;
			15'h00002E87 : data <= 8'b00000000 ;
			15'h00002E88 : data <= 8'b00000000 ;
			15'h00002E89 : data <= 8'b00000000 ;
			15'h00002E8A : data <= 8'b00000000 ;
			15'h00002E8B : data <= 8'b00000000 ;
			15'h00002E8C : data <= 8'b00000000 ;
			15'h00002E8D : data <= 8'b00000000 ;
			15'h00002E8E : data <= 8'b00000000 ;
			15'h00002E8F : data <= 8'b00000000 ;
			15'h00002E90 : data <= 8'b00000000 ;
			15'h00002E91 : data <= 8'b00000000 ;
			15'h00002E92 : data <= 8'b00000000 ;
			15'h00002E93 : data <= 8'b00000000 ;
			15'h00002E94 : data <= 8'b00000000 ;
			15'h00002E95 : data <= 8'b00000000 ;
			15'h00002E96 : data <= 8'b00000000 ;
			15'h00002E97 : data <= 8'b00000000 ;
			15'h00002E98 : data <= 8'b00000000 ;
			15'h00002E99 : data <= 8'b00000000 ;
			15'h00002E9A : data <= 8'b00000000 ;
			15'h00002E9B : data <= 8'b00000000 ;
			15'h00002E9C : data <= 8'b00000000 ;
			15'h00002E9D : data <= 8'b00000000 ;
			15'h00002E9E : data <= 8'b00000000 ;
			15'h00002E9F : data <= 8'b00000000 ;
			15'h00002EA0 : data <= 8'b00000000 ;
			15'h00002EA1 : data <= 8'b00000000 ;
			15'h00002EA2 : data <= 8'b00000000 ;
			15'h00002EA3 : data <= 8'b00000000 ;
			15'h00002EA4 : data <= 8'b00000000 ;
			15'h00002EA5 : data <= 8'b00000000 ;
			15'h00002EA6 : data <= 8'b00000000 ;
			15'h00002EA7 : data <= 8'b00000000 ;
			15'h00002EA8 : data <= 8'b00000000 ;
			15'h00002EA9 : data <= 8'b00000000 ;
			15'h00002EAA : data <= 8'b00000000 ;
			15'h00002EAB : data <= 8'b00000000 ;
			15'h00002EAC : data <= 8'b00000000 ;
			15'h00002EAD : data <= 8'b00000000 ;
			15'h00002EAE : data <= 8'b00000000 ;
			15'h00002EAF : data <= 8'b00000000 ;
			15'h00002EB0 : data <= 8'b00000000 ;
			15'h00002EB1 : data <= 8'b00000000 ;
			15'h00002EB2 : data <= 8'b00000000 ;
			15'h00002EB3 : data <= 8'b00000000 ;
			15'h00002EB4 : data <= 8'b00000000 ;
			15'h00002EB5 : data <= 8'b00000000 ;
			15'h00002EB6 : data <= 8'b00000000 ;
			15'h00002EB7 : data <= 8'b00000000 ;
			15'h00002EB8 : data <= 8'b00000000 ;
			15'h00002EB9 : data <= 8'b00000000 ;
			15'h00002EBA : data <= 8'b00000000 ;
			15'h00002EBB : data <= 8'b00000000 ;
			15'h00002EBC : data <= 8'b00000000 ;
			15'h00002EBD : data <= 8'b00000000 ;
			15'h00002EBE : data <= 8'b00000000 ;
			15'h00002EBF : data <= 8'b00000000 ;
			15'h00002EC0 : data <= 8'b00000000 ;
			15'h00002EC1 : data <= 8'b00000000 ;
			15'h00002EC2 : data <= 8'b00000000 ;
			15'h00002EC3 : data <= 8'b00000000 ;
			15'h00002EC4 : data <= 8'b00000000 ;
			15'h00002EC5 : data <= 8'b00000000 ;
			15'h00002EC6 : data <= 8'b00000000 ;
			15'h00002EC7 : data <= 8'b00000000 ;
			15'h00002EC8 : data <= 8'b00000000 ;
			15'h00002EC9 : data <= 8'b00000000 ;
			15'h00002ECA : data <= 8'b00000000 ;
			15'h00002ECB : data <= 8'b00000000 ;
			15'h00002ECC : data <= 8'b00000000 ;
			15'h00002ECD : data <= 8'b00000000 ;
			15'h00002ECE : data <= 8'b00000000 ;
			15'h00002ECF : data <= 8'b00000000 ;
			15'h00002ED0 : data <= 8'b00000000 ;
			15'h00002ED1 : data <= 8'b00000000 ;
			15'h00002ED2 : data <= 8'b00000000 ;
			15'h00002ED3 : data <= 8'b00000000 ;
			15'h00002ED4 : data <= 8'b00000000 ;
			15'h00002ED5 : data <= 8'b00000000 ;
			15'h00002ED6 : data <= 8'b00000000 ;
			15'h00002ED7 : data <= 8'b00000000 ;
			15'h00002ED8 : data <= 8'b00000000 ;
			15'h00002ED9 : data <= 8'b00000000 ;
			15'h00002EDA : data <= 8'b00000000 ;
			15'h00002EDB : data <= 8'b00000000 ;
			15'h00002EDC : data <= 8'b00000000 ;
			15'h00002EDD : data <= 8'b00000000 ;
			15'h00002EDE : data <= 8'b00000000 ;
			15'h00002EDF : data <= 8'b00000000 ;
			15'h00002EE0 : data <= 8'b00000000 ;
			15'h00002EE1 : data <= 8'b00000000 ;
			15'h00002EE2 : data <= 8'b00000000 ;
			15'h00002EE3 : data <= 8'b00000000 ;
			15'h00002EE4 : data <= 8'b00000000 ;
			15'h00002EE5 : data <= 8'b00000000 ;
			15'h00002EE6 : data <= 8'b00000000 ;
			15'h00002EE7 : data <= 8'b00000000 ;
			15'h00002EE8 : data <= 8'b00000000 ;
			15'h00002EE9 : data <= 8'b00000000 ;
			15'h00002EEA : data <= 8'b00000000 ;
			15'h00002EEB : data <= 8'b00000000 ;
			15'h00002EEC : data <= 8'b00000000 ;
			15'h00002EED : data <= 8'b00000000 ;
			15'h00002EEE : data <= 8'b00000000 ;
			15'h00002EEF : data <= 8'b00000000 ;
			15'h00002EF0 : data <= 8'b00000000 ;
			15'h00002EF1 : data <= 8'b00000000 ;
			15'h00002EF2 : data <= 8'b00000000 ;
			15'h00002EF3 : data <= 8'b00000000 ;
			15'h00002EF4 : data <= 8'b00000000 ;
			15'h00002EF5 : data <= 8'b00000000 ;
			15'h00002EF6 : data <= 8'b00000000 ;
			15'h00002EF7 : data <= 8'b00000000 ;
			15'h00002EF8 : data <= 8'b00000000 ;
			15'h00002EF9 : data <= 8'b00000000 ;
			15'h00002EFA : data <= 8'b00000000 ;
			15'h00002EFB : data <= 8'b00000000 ;
			15'h00002EFC : data <= 8'b00000000 ;
			15'h00002EFD : data <= 8'b00000000 ;
			15'h00002EFE : data <= 8'b00000000 ;
			15'h00002EFF : data <= 8'b00000000 ;
			15'h00002F00 : data <= 8'b00000000 ;
			15'h00002F01 : data <= 8'b00000000 ;
			15'h00002F02 : data <= 8'b00000000 ;
			15'h00002F03 : data <= 8'b00000000 ;
			15'h00002F04 : data <= 8'b00000000 ;
			15'h00002F05 : data <= 8'b00000000 ;
			15'h00002F06 : data <= 8'b00000000 ;
			15'h00002F07 : data <= 8'b00000000 ;
			15'h00002F08 : data <= 8'b00000000 ;
			15'h00002F09 : data <= 8'b00000000 ;
			15'h00002F0A : data <= 8'b00000000 ;
			15'h00002F0B : data <= 8'b00000000 ;
			15'h00002F0C : data <= 8'b00000000 ;
			15'h00002F0D : data <= 8'b00000000 ;
			15'h00002F0E : data <= 8'b00000000 ;
			15'h00002F0F : data <= 8'b00000000 ;
			15'h00002F10 : data <= 8'b00000000 ;
			15'h00002F11 : data <= 8'b00000000 ;
			15'h00002F12 : data <= 8'b00000000 ;
			15'h00002F13 : data <= 8'b00000000 ;
			15'h00002F14 : data <= 8'b00000000 ;
			15'h00002F15 : data <= 8'b00000000 ;
			15'h00002F16 : data <= 8'b00000000 ;
			15'h00002F17 : data <= 8'b00000000 ;
			15'h00002F18 : data <= 8'b00000000 ;
			15'h00002F19 : data <= 8'b00000000 ;
			15'h00002F1A : data <= 8'b00000000 ;
			15'h00002F1B : data <= 8'b00000000 ;
			15'h00002F1C : data <= 8'b00000000 ;
			15'h00002F1D : data <= 8'b00000000 ;
			15'h00002F1E : data <= 8'b00000000 ;
			15'h00002F1F : data <= 8'b00000000 ;
			15'h00002F20 : data <= 8'b00000000 ;
			15'h00002F21 : data <= 8'b00000000 ;
			15'h00002F22 : data <= 8'b00000000 ;
			15'h00002F23 : data <= 8'b00000000 ;
			15'h00002F24 : data <= 8'b00000000 ;
			15'h00002F25 : data <= 8'b00000000 ;
			15'h00002F26 : data <= 8'b00000000 ;
			15'h00002F27 : data <= 8'b00000000 ;
			15'h00002F28 : data <= 8'b00000000 ;
			15'h00002F29 : data <= 8'b00000000 ;
			15'h00002F2A : data <= 8'b00000000 ;
			15'h00002F2B : data <= 8'b00000000 ;
			15'h00002F2C : data <= 8'b00000000 ;
			15'h00002F2D : data <= 8'b00000000 ;
			15'h00002F2E : data <= 8'b00000000 ;
			15'h00002F2F : data <= 8'b00000000 ;
			15'h00002F30 : data <= 8'b00000000 ;
			15'h00002F31 : data <= 8'b00000000 ;
			15'h00002F32 : data <= 8'b00000000 ;
			15'h00002F33 : data <= 8'b00000000 ;
			15'h00002F34 : data <= 8'b00000000 ;
			15'h00002F35 : data <= 8'b00000000 ;
			15'h00002F36 : data <= 8'b00000000 ;
			15'h00002F37 : data <= 8'b00000000 ;
			15'h00002F38 : data <= 8'b00000000 ;
			15'h00002F39 : data <= 8'b00000000 ;
			15'h00002F3A : data <= 8'b00000000 ;
			15'h00002F3B : data <= 8'b00000000 ;
			15'h00002F3C : data <= 8'b00000000 ;
			15'h00002F3D : data <= 8'b00000000 ;
			15'h00002F3E : data <= 8'b00000000 ;
			15'h00002F3F : data <= 8'b00000000 ;
			15'h00002F40 : data <= 8'b00000000 ;
			15'h00002F41 : data <= 8'b00000000 ;
			15'h00002F42 : data <= 8'b00000000 ;
			15'h00002F43 : data <= 8'b00000000 ;
			15'h00002F44 : data <= 8'b00000000 ;
			15'h00002F45 : data <= 8'b00000000 ;
			15'h00002F46 : data <= 8'b00000000 ;
			15'h00002F47 : data <= 8'b00000000 ;
			15'h00002F48 : data <= 8'b00000000 ;
			15'h00002F49 : data <= 8'b00000000 ;
			15'h00002F4A : data <= 8'b00000000 ;
			15'h00002F4B : data <= 8'b00000000 ;
			15'h00002F4C : data <= 8'b00000000 ;
			15'h00002F4D : data <= 8'b00000000 ;
			15'h00002F4E : data <= 8'b00000000 ;
			15'h00002F4F : data <= 8'b00000000 ;
			15'h00002F50 : data <= 8'b00000000 ;
			15'h00002F51 : data <= 8'b00000000 ;
			15'h00002F52 : data <= 8'b00000000 ;
			15'h00002F53 : data <= 8'b00000000 ;
			15'h00002F54 : data <= 8'b00000000 ;
			15'h00002F55 : data <= 8'b00000000 ;
			15'h00002F56 : data <= 8'b00000000 ;
			15'h00002F57 : data <= 8'b00000000 ;
			15'h00002F58 : data <= 8'b00000000 ;
			15'h00002F59 : data <= 8'b00000000 ;
			15'h00002F5A : data <= 8'b00000000 ;
			15'h00002F5B : data <= 8'b00000000 ;
			15'h00002F5C : data <= 8'b00000000 ;
			15'h00002F5D : data <= 8'b00000000 ;
			15'h00002F5E : data <= 8'b00000000 ;
			15'h00002F5F : data <= 8'b00000000 ;
			15'h00002F60 : data <= 8'b00000000 ;
			15'h00002F61 : data <= 8'b00000000 ;
			15'h00002F62 : data <= 8'b00000000 ;
			15'h00002F63 : data <= 8'b00000000 ;
			15'h00002F64 : data <= 8'b00000000 ;
			15'h00002F65 : data <= 8'b00000000 ;
			15'h00002F66 : data <= 8'b00000000 ;
			15'h00002F67 : data <= 8'b00000000 ;
			15'h00002F68 : data <= 8'b00000000 ;
			15'h00002F69 : data <= 8'b00000000 ;
			15'h00002F6A : data <= 8'b00000000 ;
			15'h00002F6B : data <= 8'b00000000 ;
			15'h00002F6C : data <= 8'b00000000 ;
			15'h00002F6D : data <= 8'b00000000 ;
			15'h00002F6E : data <= 8'b00000000 ;
			15'h00002F6F : data <= 8'b00000000 ;
			15'h00002F70 : data <= 8'b00000000 ;
			15'h00002F71 : data <= 8'b00000000 ;
			15'h00002F72 : data <= 8'b00000000 ;
			15'h00002F73 : data <= 8'b00000000 ;
			15'h00002F74 : data <= 8'b00000000 ;
			15'h00002F75 : data <= 8'b00000000 ;
			15'h00002F76 : data <= 8'b00000000 ;
			15'h00002F77 : data <= 8'b00000000 ;
			15'h00002F78 : data <= 8'b00000000 ;
			15'h00002F79 : data <= 8'b00000000 ;
			15'h00002F7A : data <= 8'b00000000 ;
			15'h00002F7B : data <= 8'b00000000 ;
			15'h00002F7C : data <= 8'b00000000 ;
			15'h00002F7D : data <= 8'b00000000 ;
			15'h00002F7E : data <= 8'b00000000 ;
			15'h00002F7F : data <= 8'b00000000 ;
			15'h00002F80 : data <= 8'b00000000 ;
			15'h00002F81 : data <= 8'b00000000 ;
			15'h00002F82 : data <= 8'b00000000 ;
			15'h00002F83 : data <= 8'b00000000 ;
			15'h00002F84 : data <= 8'b00000000 ;
			15'h00002F85 : data <= 8'b00000000 ;
			15'h00002F86 : data <= 8'b00000000 ;
			15'h00002F87 : data <= 8'b00000000 ;
			15'h00002F88 : data <= 8'b00000000 ;
			15'h00002F89 : data <= 8'b00000000 ;
			15'h00002F8A : data <= 8'b00000000 ;
			15'h00002F8B : data <= 8'b00000000 ;
			15'h00002F8C : data <= 8'b00000000 ;
			15'h00002F8D : data <= 8'b00000000 ;
			15'h00002F8E : data <= 8'b00000000 ;
			15'h00002F8F : data <= 8'b00000000 ;
			15'h00002F90 : data <= 8'b00000000 ;
			15'h00002F91 : data <= 8'b00000000 ;
			15'h00002F92 : data <= 8'b00000000 ;
			15'h00002F93 : data <= 8'b00000000 ;
			15'h00002F94 : data <= 8'b00000000 ;
			15'h00002F95 : data <= 8'b00000000 ;
			15'h00002F96 : data <= 8'b00000000 ;
			15'h00002F97 : data <= 8'b00000000 ;
			15'h00002F98 : data <= 8'b00000000 ;
			15'h00002F99 : data <= 8'b00000000 ;
			15'h00002F9A : data <= 8'b00000000 ;
			15'h00002F9B : data <= 8'b00000000 ;
			15'h00002F9C : data <= 8'b00000000 ;
			15'h00002F9D : data <= 8'b00000000 ;
			15'h00002F9E : data <= 8'b00000000 ;
			15'h00002F9F : data <= 8'b00000000 ;
			15'h00002FA0 : data <= 8'b00000000 ;
			15'h00002FA1 : data <= 8'b00000000 ;
			15'h00002FA2 : data <= 8'b00000000 ;
			15'h00002FA3 : data <= 8'b00000000 ;
			15'h00002FA4 : data <= 8'b00000000 ;
			15'h00002FA5 : data <= 8'b00000000 ;
			15'h00002FA6 : data <= 8'b00000000 ;
			15'h00002FA7 : data <= 8'b00000000 ;
			15'h00002FA8 : data <= 8'b00000000 ;
			15'h00002FA9 : data <= 8'b00000000 ;
			15'h00002FAA : data <= 8'b00000000 ;
			15'h00002FAB : data <= 8'b00000000 ;
			15'h00002FAC : data <= 8'b00000000 ;
			15'h00002FAD : data <= 8'b00000000 ;
			15'h00002FAE : data <= 8'b00000000 ;
			15'h00002FAF : data <= 8'b00000000 ;
			15'h00002FB0 : data <= 8'b00000000 ;
			15'h00002FB1 : data <= 8'b00000000 ;
			15'h00002FB2 : data <= 8'b00000000 ;
			15'h00002FB3 : data <= 8'b00000000 ;
			15'h00002FB4 : data <= 8'b00000000 ;
			15'h00002FB5 : data <= 8'b00000000 ;
			15'h00002FB6 : data <= 8'b00000000 ;
			15'h00002FB7 : data <= 8'b00000000 ;
			15'h00002FB8 : data <= 8'b00000000 ;
			15'h00002FB9 : data <= 8'b00000000 ;
			15'h00002FBA : data <= 8'b00000000 ;
			15'h00002FBB : data <= 8'b00000000 ;
			15'h00002FBC : data <= 8'b00000000 ;
			15'h00002FBD : data <= 8'b00000000 ;
			15'h00002FBE : data <= 8'b00000000 ;
			15'h00002FBF : data <= 8'b00000000 ;
			15'h00002FC0 : data <= 8'b00000000 ;
			15'h00002FC1 : data <= 8'b00000000 ;
			15'h00002FC2 : data <= 8'b00000000 ;
			15'h00002FC3 : data <= 8'b00000000 ;
			15'h00002FC4 : data <= 8'b00000000 ;
			15'h00002FC5 : data <= 8'b00000000 ;
			15'h00002FC6 : data <= 8'b00000000 ;
			15'h00002FC7 : data <= 8'b00000000 ;
			15'h00002FC8 : data <= 8'b00000000 ;
			15'h00002FC9 : data <= 8'b00000000 ;
			15'h00002FCA : data <= 8'b00000000 ;
			15'h00002FCB : data <= 8'b00000000 ;
			15'h00002FCC : data <= 8'b00000000 ;
			15'h00002FCD : data <= 8'b00000000 ;
			15'h00002FCE : data <= 8'b00000000 ;
			15'h00002FCF : data <= 8'b00000000 ;
			15'h00002FD0 : data <= 8'b00000000 ;
			15'h00002FD1 : data <= 8'b00000000 ;
			15'h00002FD2 : data <= 8'b00000000 ;
			15'h00002FD3 : data <= 8'b00000000 ;
			15'h00002FD4 : data <= 8'b00000000 ;
			15'h00002FD5 : data <= 8'b00000000 ;
			15'h00002FD6 : data <= 8'b00000000 ;
			15'h00002FD7 : data <= 8'b00000000 ;
			15'h00002FD8 : data <= 8'b00000000 ;
			15'h00002FD9 : data <= 8'b00000000 ;
			15'h00002FDA : data <= 8'b00000000 ;
			15'h00002FDB : data <= 8'b00000000 ;
			15'h00002FDC : data <= 8'b00000000 ;
			15'h00002FDD : data <= 8'b00000000 ;
			15'h00002FDE : data <= 8'b00000000 ;
			15'h00002FDF : data <= 8'b00000000 ;
			15'h00002FE0 : data <= 8'b00000000 ;
			15'h00002FE1 : data <= 8'b00000000 ;
			15'h00002FE2 : data <= 8'b00000000 ;
			15'h00002FE3 : data <= 8'b00000000 ;
			15'h00002FE4 : data <= 8'b00000000 ;
			15'h00002FE5 : data <= 8'b00000000 ;
			15'h00002FE6 : data <= 8'b00000000 ;
			15'h00002FE7 : data <= 8'b00000000 ;
			15'h00002FE8 : data <= 8'b00000000 ;
			15'h00002FE9 : data <= 8'b00000000 ;
			15'h00002FEA : data <= 8'b00000000 ;
			15'h00002FEB : data <= 8'b00000000 ;
			15'h00002FEC : data <= 8'b00000000 ;
			15'h00002FED : data <= 8'b00000000 ;
			15'h00002FEE : data <= 8'b00000000 ;
			15'h00002FEF : data <= 8'b00000000 ;
			15'h00002FF0 : data <= 8'b00000000 ;
			15'h00002FF1 : data <= 8'b00000000 ;
			15'h00002FF2 : data <= 8'b00000000 ;
			15'h00002FF3 : data <= 8'b00000000 ;
			15'h00002FF4 : data <= 8'b00000000 ;
			15'h00002FF5 : data <= 8'b00000000 ;
			15'h00002FF6 : data <= 8'b00000000 ;
			15'h00002FF7 : data <= 8'b00000000 ;
			15'h00002FF8 : data <= 8'b00000000 ;
			15'h00002FF9 : data <= 8'b00000000 ;
			15'h00002FFA : data <= 8'b00000000 ;
			15'h00002FFB : data <= 8'b00000000 ;
			15'h00002FFC : data <= 8'b00000000 ;
			15'h00002FFD : data <= 8'b00000000 ;
			15'h00002FFE : data <= 8'b00000000 ;
			15'h00002FFF : data <= 8'b00000000 ;
			15'h00003000 : data <= 8'b00000000 ;
			15'h00003001 : data <= 8'b00000000 ;
			15'h00003002 : data <= 8'b00000000 ;
			15'h00003003 : data <= 8'b00000000 ;
			15'h00003004 : data <= 8'b00000000 ;
			15'h00003005 : data <= 8'b00000000 ;
			15'h00003006 : data <= 8'b00000000 ;
			15'h00003007 : data <= 8'b00000000 ;
			15'h00003008 : data <= 8'b00000000 ;
			15'h00003009 : data <= 8'b00000000 ;
			15'h0000300A : data <= 8'b00000000 ;
			15'h0000300B : data <= 8'b00000000 ;
			15'h0000300C : data <= 8'b00000000 ;
			15'h0000300D : data <= 8'b00000000 ;
			15'h0000300E : data <= 8'b00000000 ;
			15'h0000300F : data <= 8'b00000000 ;
			15'h00003010 : data <= 8'b00000000 ;
			15'h00003011 : data <= 8'b00000000 ;
			15'h00003012 : data <= 8'b00000000 ;
			15'h00003013 : data <= 8'b00000000 ;
			15'h00003014 : data <= 8'b00000000 ;
			15'h00003015 : data <= 8'b00000000 ;
			15'h00003016 : data <= 8'b00000000 ;
			15'h00003017 : data <= 8'b00000000 ;
			15'h00003018 : data <= 8'b00000000 ;
			15'h00003019 : data <= 8'b00000000 ;
			15'h0000301A : data <= 8'b00000000 ;
			15'h0000301B : data <= 8'b00000000 ;
			15'h0000301C : data <= 8'b00000000 ;
			15'h0000301D : data <= 8'b00000000 ;
			15'h0000301E : data <= 8'b00000000 ;
			15'h0000301F : data <= 8'b00000000 ;
			15'h00003020 : data <= 8'b00000000 ;
			15'h00003021 : data <= 8'b00000000 ;
			15'h00003022 : data <= 8'b00000000 ;
			15'h00003023 : data <= 8'b00000000 ;
			15'h00003024 : data <= 8'b00000000 ;
			15'h00003025 : data <= 8'b00000000 ;
			15'h00003026 : data <= 8'b00000000 ;
			15'h00003027 : data <= 8'b00000000 ;
			15'h00003028 : data <= 8'b00000000 ;
			15'h00003029 : data <= 8'b00000000 ;
			15'h0000302A : data <= 8'b00000000 ;
			15'h0000302B : data <= 8'b00000000 ;
			15'h0000302C : data <= 8'b00000000 ;
			15'h0000302D : data <= 8'b00000000 ;
			15'h0000302E : data <= 8'b00000000 ;
			15'h0000302F : data <= 8'b00000000 ;
			15'h00003030 : data <= 8'b00000000 ;
			15'h00003031 : data <= 8'b00000000 ;
			15'h00003032 : data <= 8'b00000000 ;
			15'h00003033 : data <= 8'b00000000 ;
			15'h00003034 : data <= 8'b00000000 ;
			15'h00003035 : data <= 8'b00000000 ;
			15'h00003036 : data <= 8'b00000000 ;
			15'h00003037 : data <= 8'b00000000 ;
			15'h00003038 : data <= 8'b00000000 ;
			15'h00003039 : data <= 8'b00000000 ;
			15'h0000303A : data <= 8'b00000000 ;
			15'h0000303B : data <= 8'b00000000 ;
			15'h0000303C : data <= 8'b00000000 ;
			15'h0000303D : data <= 8'b00000000 ;
			15'h0000303E : data <= 8'b00000000 ;
			15'h0000303F : data <= 8'b00000000 ;
			15'h00003040 : data <= 8'b00000000 ;
			15'h00003041 : data <= 8'b00000000 ;
			15'h00003042 : data <= 8'b00000000 ;
			15'h00003043 : data <= 8'b00000000 ;
			15'h00003044 : data <= 8'b00000000 ;
			15'h00003045 : data <= 8'b00000000 ;
			15'h00003046 : data <= 8'b00000000 ;
			15'h00003047 : data <= 8'b00000000 ;
			15'h00003048 : data <= 8'b00000000 ;
			15'h00003049 : data <= 8'b00000000 ;
			15'h0000304A : data <= 8'b00000000 ;
			15'h0000304B : data <= 8'b00000000 ;
			15'h0000304C : data <= 8'b00000000 ;
			15'h0000304D : data <= 8'b00000000 ;
			15'h0000304E : data <= 8'b00000000 ;
			15'h0000304F : data <= 8'b00000000 ;
			15'h00003050 : data <= 8'b00000000 ;
			15'h00003051 : data <= 8'b00000000 ;
			15'h00003052 : data <= 8'b00000000 ;
			15'h00003053 : data <= 8'b00000000 ;
			15'h00003054 : data <= 8'b00000000 ;
			15'h00003055 : data <= 8'b00000000 ;
			15'h00003056 : data <= 8'b00000000 ;
			15'h00003057 : data <= 8'b00000000 ;
			15'h00003058 : data <= 8'b00000000 ;
			15'h00003059 : data <= 8'b00000000 ;
			15'h0000305A : data <= 8'b00000000 ;
			15'h0000305B : data <= 8'b00000000 ;
			15'h0000305C : data <= 8'b00000000 ;
			15'h0000305D : data <= 8'b00000000 ;
			15'h0000305E : data <= 8'b00000000 ;
			15'h0000305F : data <= 8'b00000000 ;
			15'h00003060 : data <= 8'b00000000 ;
			15'h00003061 : data <= 8'b00000000 ;
			15'h00003062 : data <= 8'b00000000 ;
			15'h00003063 : data <= 8'b00000000 ;
			15'h00003064 : data <= 8'b00000000 ;
			15'h00003065 : data <= 8'b00000000 ;
			15'h00003066 : data <= 8'b00000000 ;
			15'h00003067 : data <= 8'b00000000 ;
			15'h00003068 : data <= 8'b00000000 ;
			15'h00003069 : data <= 8'b00000000 ;
			15'h0000306A : data <= 8'b00000000 ;
			15'h0000306B : data <= 8'b00000000 ;
			15'h0000306C : data <= 8'b00000000 ;
			15'h0000306D : data <= 8'b00000000 ;
			15'h0000306E : data <= 8'b00000000 ;
			15'h0000306F : data <= 8'b00000000 ;
			15'h00003070 : data <= 8'b00000000 ;
			15'h00003071 : data <= 8'b00000000 ;
			15'h00003072 : data <= 8'b00000000 ;
			15'h00003073 : data <= 8'b00000000 ;
			15'h00003074 : data <= 8'b00000000 ;
			15'h00003075 : data <= 8'b00000000 ;
			15'h00003076 : data <= 8'b00000000 ;
			15'h00003077 : data <= 8'b00000000 ;
			15'h00003078 : data <= 8'b00000000 ;
			15'h00003079 : data <= 8'b00000000 ;
			15'h0000307A : data <= 8'b00000000 ;
			15'h0000307B : data <= 8'b00000000 ;
			15'h0000307C : data <= 8'b00000000 ;
			15'h0000307D : data <= 8'b00000000 ;
			15'h0000307E : data <= 8'b00000000 ;
			15'h0000307F : data <= 8'b00000000 ;
			15'h00003080 : data <= 8'b00000000 ;
			15'h00003081 : data <= 8'b00000000 ;
			15'h00003082 : data <= 8'b00000000 ;
			15'h00003083 : data <= 8'b00000000 ;
			15'h00003084 : data <= 8'b00000000 ;
			15'h00003085 : data <= 8'b00000000 ;
			15'h00003086 : data <= 8'b00000000 ;
			15'h00003087 : data <= 8'b00000000 ;
			15'h00003088 : data <= 8'b00000000 ;
			15'h00003089 : data <= 8'b00000000 ;
			15'h0000308A : data <= 8'b00000000 ;
			15'h0000308B : data <= 8'b00000000 ;
			15'h0000308C : data <= 8'b00000000 ;
			15'h0000308D : data <= 8'b00000000 ;
			15'h0000308E : data <= 8'b00000000 ;
			15'h0000308F : data <= 8'b00000000 ;
			15'h00003090 : data <= 8'b00000000 ;
			15'h00003091 : data <= 8'b00000000 ;
			15'h00003092 : data <= 8'b00000000 ;
			15'h00003093 : data <= 8'b00000000 ;
			15'h00003094 : data <= 8'b00000000 ;
			15'h00003095 : data <= 8'b00000000 ;
			15'h00003096 : data <= 8'b00000000 ;
			15'h00003097 : data <= 8'b00000000 ;
			15'h00003098 : data <= 8'b00000000 ;
			15'h00003099 : data <= 8'b00000000 ;
			15'h0000309A : data <= 8'b00000000 ;
			15'h0000309B : data <= 8'b00000000 ;
			15'h0000309C : data <= 8'b00000000 ;
			15'h0000309D : data <= 8'b00000000 ;
			15'h0000309E : data <= 8'b00000000 ;
			15'h0000309F : data <= 8'b00000000 ;
			15'h000030A0 : data <= 8'b00000000 ;
			15'h000030A1 : data <= 8'b00000000 ;
			15'h000030A2 : data <= 8'b00000000 ;
			15'h000030A3 : data <= 8'b00000000 ;
			15'h000030A4 : data <= 8'b00000000 ;
			15'h000030A5 : data <= 8'b00000000 ;
			15'h000030A6 : data <= 8'b00000000 ;
			15'h000030A7 : data <= 8'b00000000 ;
			15'h000030A8 : data <= 8'b00000000 ;
			15'h000030A9 : data <= 8'b00000000 ;
			15'h000030AA : data <= 8'b00000000 ;
			15'h000030AB : data <= 8'b00000000 ;
			15'h000030AC : data <= 8'b00000000 ;
			15'h000030AD : data <= 8'b00000000 ;
			15'h000030AE : data <= 8'b00000000 ;
			15'h000030AF : data <= 8'b00000000 ;
			15'h000030B0 : data <= 8'b00000000 ;
			15'h000030B1 : data <= 8'b00000000 ;
			15'h000030B2 : data <= 8'b00000000 ;
			15'h000030B3 : data <= 8'b00000000 ;
			15'h000030B4 : data <= 8'b00000000 ;
			15'h000030B5 : data <= 8'b00000000 ;
			15'h000030B6 : data <= 8'b00000000 ;
			15'h000030B7 : data <= 8'b00000000 ;
			15'h000030B8 : data <= 8'b00000000 ;
			15'h000030B9 : data <= 8'b00000000 ;
			15'h000030BA : data <= 8'b00000000 ;
			15'h000030BB : data <= 8'b00000000 ;
			15'h000030BC : data <= 8'b00000000 ;
			15'h000030BD : data <= 8'b00000000 ;
			15'h000030BE : data <= 8'b00000000 ;
			15'h000030BF : data <= 8'b00000000 ;
			15'h000030C0 : data <= 8'b00000000 ;
			15'h000030C1 : data <= 8'b00000000 ;
			15'h000030C2 : data <= 8'b00000000 ;
			15'h000030C3 : data <= 8'b00000000 ;
			15'h000030C4 : data <= 8'b00000000 ;
			15'h000030C5 : data <= 8'b00000000 ;
			15'h000030C6 : data <= 8'b00000000 ;
			15'h000030C7 : data <= 8'b00000000 ;
			15'h000030C8 : data <= 8'b00000000 ;
			15'h000030C9 : data <= 8'b00000000 ;
			15'h000030CA : data <= 8'b00000000 ;
			15'h000030CB : data <= 8'b00000000 ;
			15'h000030CC : data <= 8'b00000000 ;
			15'h000030CD : data <= 8'b00000000 ;
			15'h000030CE : data <= 8'b00000000 ;
			15'h000030CF : data <= 8'b00000000 ;
			15'h000030D0 : data <= 8'b00000000 ;
			15'h000030D1 : data <= 8'b00000000 ;
			15'h000030D2 : data <= 8'b00000000 ;
			15'h000030D3 : data <= 8'b00000000 ;
			15'h000030D4 : data <= 8'b00000000 ;
			15'h000030D5 : data <= 8'b00000000 ;
			15'h000030D6 : data <= 8'b00000000 ;
			15'h000030D7 : data <= 8'b00000000 ;
			15'h000030D8 : data <= 8'b00000000 ;
			15'h000030D9 : data <= 8'b00000000 ;
			15'h000030DA : data <= 8'b00000000 ;
			15'h000030DB : data <= 8'b00000000 ;
			15'h000030DC : data <= 8'b00000000 ;
			15'h000030DD : data <= 8'b00000000 ;
			15'h000030DE : data <= 8'b00000000 ;
			15'h000030DF : data <= 8'b00000000 ;
			15'h000030E0 : data <= 8'b00000000 ;
			15'h000030E1 : data <= 8'b00000000 ;
			15'h000030E2 : data <= 8'b00000000 ;
			15'h000030E3 : data <= 8'b00000000 ;
			15'h000030E4 : data <= 8'b00000000 ;
			15'h000030E5 : data <= 8'b00000000 ;
			15'h000030E6 : data <= 8'b00000000 ;
			15'h000030E7 : data <= 8'b00000000 ;
			15'h000030E8 : data <= 8'b00000000 ;
			15'h000030E9 : data <= 8'b00000000 ;
			15'h000030EA : data <= 8'b00000000 ;
			15'h000030EB : data <= 8'b00000000 ;
			15'h000030EC : data <= 8'b00000000 ;
			15'h000030ED : data <= 8'b00000000 ;
			15'h000030EE : data <= 8'b00000000 ;
			15'h000030EF : data <= 8'b00000000 ;
			15'h000030F0 : data <= 8'b00000000 ;
			15'h000030F1 : data <= 8'b00000000 ;
			15'h000030F2 : data <= 8'b00000000 ;
			15'h000030F3 : data <= 8'b00000000 ;
			15'h000030F4 : data <= 8'b00000000 ;
			15'h000030F5 : data <= 8'b00000000 ;
			15'h000030F6 : data <= 8'b00000000 ;
			15'h000030F7 : data <= 8'b00000000 ;
			15'h000030F8 : data <= 8'b00000000 ;
			15'h000030F9 : data <= 8'b00000000 ;
			15'h000030FA : data <= 8'b00000000 ;
			15'h000030FB : data <= 8'b00000000 ;
			15'h000030FC : data <= 8'b00000000 ;
			15'h000030FD : data <= 8'b00000000 ;
			15'h000030FE : data <= 8'b00000000 ;
			15'h000030FF : data <= 8'b00000000 ;
			15'h00003100 : data <= 8'b00000000 ;
			15'h00003101 : data <= 8'b00000000 ;
			15'h00003102 : data <= 8'b00000000 ;
			15'h00003103 : data <= 8'b00000000 ;
			15'h00003104 : data <= 8'b00000000 ;
			15'h00003105 : data <= 8'b00000000 ;
			15'h00003106 : data <= 8'b00000000 ;
			15'h00003107 : data <= 8'b00000000 ;
			15'h00003108 : data <= 8'b00000000 ;
			15'h00003109 : data <= 8'b00000000 ;
			15'h0000310A : data <= 8'b00000000 ;
			15'h0000310B : data <= 8'b00000000 ;
			15'h0000310C : data <= 8'b00000000 ;
			15'h0000310D : data <= 8'b00000000 ;
			15'h0000310E : data <= 8'b00000000 ;
			15'h0000310F : data <= 8'b00000000 ;
			15'h00003110 : data <= 8'b00000000 ;
			15'h00003111 : data <= 8'b00000000 ;
			15'h00003112 : data <= 8'b00000000 ;
			15'h00003113 : data <= 8'b00000000 ;
			15'h00003114 : data <= 8'b00000000 ;
			15'h00003115 : data <= 8'b00000000 ;
			15'h00003116 : data <= 8'b00000000 ;
			15'h00003117 : data <= 8'b00000000 ;
			15'h00003118 : data <= 8'b00000000 ;
			15'h00003119 : data <= 8'b00000000 ;
			15'h0000311A : data <= 8'b00000000 ;
			15'h0000311B : data <= 8'b00000000 ;
			15'h0000311C : data <= 8'b00000000 ;
			15'h0000311D : data <= 8'b00000000 ;
			15'h0000311E : data <= 8'b00000000 ;
			15'h0000311F : data <= 8'b00000000 ;
			15'h00003120 : data <= 8'b00000000 ;
			15'h00003121 : data <= 8'b00000000 ;
			15'h00003122 : data <= 8'b00000000 ;
			15'h00003123 : data <= 8'b00000000 ;
			15'h00003124 : data <= 8'b00000000 ;
			15'h00003125 : data <= 8'b00000000 ;
			15'h00003126 : data <= 8'b00000000 ;
			15'h00003127 : data <= 8'b00000000 ;
			15'h00003128 : data <= 8'b00000000 ;
			15'h00003129 : data <= 8'b00000000 ;
			15'h0000312A : data <= 8'b00000000 ;
			15'h0000312B : data <= 8'b00000000 ;
			15'h0000312C : data <= 8'b00000000 ;
			15'h0000312D : data <= 8'b00000000 ;
			15'h0000312E : data <= 8'b00000000 ;
			15'h0000312F : data <= 8'b00000000 ;
			15'h00003130 : data <= 8'b00000000 ;
			15'h00003131 : data <= 8'b00000000 ;
			15'h00003132 : data <= 8'b00000000 ;
			15'h00003133 : data <= 8'b00000000 ;
			15'h00003134 : data <= 8'b00000000 ;
			15'h00003135 : data <= 8'b00000000 ;
			15'h00003136 : data <= 8'b00000000 ;
			15'h00003137 : data <= 8'b00000000 ;
			15'h00003138 : data <= 8'b00000000 ;
			15'h00003139 : data <= 8'b00000000 ;
			15'h0000313A : data <= 8'b00000000 ;
			15'h0000313B : data <= 8'b00000000 ;
			15'h0000313C : data <= 8'b00000000 ;
			15'h0000313D : data <= 8'b00000000 ;
			15'h0000313E : data <= 8'b00000000 ;
			15'h0000313F : data <= 8'b00000000 ;
			15'h00003140 : data <= 8'b00000000 ;
			15'h00003141 : data <= 8'b00000000 ;
			15'h00003142 : data <= 8'b00000000 ;
			15'h00003143 : data <= 8'b00000000 ;
			15'h00003144 : data <= 8'b00000000 ;
			15'h00003145 : data <= 8'b00000000 ;
			15'h00003146 : data <= 8'b00000000 ;
			15'h00003147 : data <= 8'b00000000 ;
			15'h00003148 : data <= 8'b00000000 ;
			15'h00003149 : data <= 8'b00000000 ;
			15'h0000314A : data <= 8'b00000000 ;
			15'h0000314B : data <= 8'b00000000 ;
			15'h0000314C : data <= 8'b00000000 ;
			15'h0000314D : data <= 8'b00000000 ;
			15'h0000314E : data <= 8'b00000000 ;
			15'h0000314F : data <= 8'b00000000 ;
			15'h00003150 : data <= 8'b00000000 ;
			15'h00003151 : data <= 8'b00000000 ;
			15'h00003152 : data <= 8'b00000000 ;
			15'h00003153 : data <= 8'b00000000 ;
			15'h00003154 : data <= 8'b00000000 ;
			15'h00003155 : data <= 8'b00000000 ;
			15'h00003156 : data <= 8'b00000000 ;
			15'h00003157 : data <= 8'b00000000 ;
			15'h00003158 : data <= 8'b00000000 ;
			15'h00003159 : data <= 8'b00000000 ;
			15'h0000315A : data <= 8'b00000000 ;
			15'h0000315B : data <= 8'b00000000 ;
			15'h0000315C : data <= 8'b00000000 ;
			15'h0000315D : data <= 8'b00000000 ;
			15'h0000315E : data <= 8'b00000000 ;
			15'h0000315F : data <= 8'b00000000 ;
			15'h00003160 : data <= 8'b00000000 ;
			15'h00003161 : data <= 8'b00000000 ;
			15'h00003162 : data <= 8'b00000000 ;
			15'h00003163 : data <= 8'b00000000 ;
			15'h00003164 : data <= 8'b00000000 ;
			15'h00003165 : data <= 8'b00000000 ;
			15'h00003166 : data <= 8'b00000000 ;
			15'h00003167 : data <= 8'b00000000 ;
			15'h00003168 : data <= 8'b00000000 ;
			15'h00003169 : data <= 8'b00000000 ;
			15'h0000316A : data <= 8'b00000000 ;
			15'h0000316B : data <= 8'b00000000 ;
			15'h0000316C : data <= 8'b00000000 ;
			15'h0000316D : data <= 8'b00000000 ;
			15'h0000316E : data <= 8'b00000000 ;
			15'h0000316F : data <= 8'b00000000 ;
			15'h00003170 : data <= 8'b00000000 ;
			15'h00003171 : data <= 8'b00000000 ;
			15'h00003172 : data <= 8'b00000000 ;
			15'h00003173 : data <= 8'b00000000 ;
			15'h00003174 : data <= 8'b00000000 ;
			15'h00003175 : data <= 8'b00000000 ;
			15'h00003176 : data <= 8'b00000000 ;
			15'h00003177 : data <= 8'b00000000 ;
			15'h00003178 : data <= 8'b00000000 ;
			15'h00003179 : data <= 8'b00000000 ;
			15'h0000317A : data <= 8'b00000000 ;
			15'h0000317B : data <= 8'b00000000 ;
			15'h0000317C : data <= 8'b00000000 ;
			15'h0000317D : data <= 8'b00000000 ;
			15'h0000317E : data <= 8'b00000000 ;
			15'h0000317F : data <= 8'b00000000 ;
			15'h00003180 : data <= 8'b00000000 ;
			15'h00003181 : data <= 8'b00000000 ;
			15'h00003182 : data <= 8'b00000000 ;
			15'h00003183 : data <= 8'b00000000 ;
			15'h00003184 : data <= 8'b00000000 ;
			15'h00003185 : data <= 8'b00000000 ;
			15'h00003186 : data <= 8'b00000000 ;
			15'h00003187 : data <= 8'b00000000 ;
			15'h00003188 : data <= 8'b00000000 ;
			15'h00003189 : data <= 8'b00000000 ;
			15'h0000318A : data <= 8'b00000000 ;
			15'h0000318B : data <= 8'b00000000 ;
			15'h0000318C : data <= 8'b00000000 ;
			15'h0000318D : data <= 8'b00000000 ;
			15'h0000318E : data <= 8'b00000000 ;
			15'h0000318F : data <= 8'b00000000 ;
			15'h00003190 : data <= 8'b00000000 ;
			15'h00003191 : data <= 8'b00000000 ;
			15'h00003192 : data <= 8'b00000000 ;
			15'h00003193 : data <= 8'b00000000 ;
			15'h00003194 : data <= 8'b00000000 ;
			15'h00003195 : data <= 8'b00000000 ;
			15'h00003196 : data <= 8'b00000000 ;
			15'h00003197 : data <= 8'b00000000 ;
			15'h00003198 : data <= 8'b00000000 ;
			15'h00003199 : data <= 8'b00000000 ;
			15'h0000319A : data <= 8'b00000000 ;
			15'h0000319B : data <= 8'b00000000 ;
			15'h0000319C : data <= 8'b00000000 ;
			15'h0000319D : data <= 8'b00000000 ;
			15'h0000319E : data <= 8'b00000000 ;
			15'h0000319F : data <= 8'b00000000 ;
			15'h000031A0 : data <= 8'b00000000 ;
			15'h000031A1 : data <= 8'b00000000 ;
			15'h000031A2 : data <= 8'b00000000 ;
			15'h000031A3 : data <= 8'b00000000 ;
			15'h000031A4 : data <= 8'b00000000 ;
			15'h000031A5 : data <= 8'b00000000 ;
			15'h000031A6 : data <= 8'b00000000 ;
			15'h000031A7 : data <= 8'b00000000 ;
			15'h000031A8 : data <= 8'b00000000 ;
			15'h000031A9 : data <= 8'b00000000 ;
			15'h000031AA : data <= 8'b00000000 ;
			15'h000031AB : data <= 8'b00000000 ;
			15'h000031AC : data <= 8'b00000000 ;
			15'h000031AD : data <= 8'b00000000 ;
			15'h000031AE : data <= 8'b00000000 ;
			15'h000031AF : data <= 8'b00000000 ;
			15'h000031B0 : data <= 8'b00000000 ;
			15'h000031B1 : data <= 8'b00000000 ;
			15'h000031B2 : data <= 8'b00000000 ;
			15'h000031B3 : data <= 8'b00000000 ;
			15'h000031B4 : data <= 8'b00000000 ;
			15'h000031B5 : data <= 8'b00000000 ;
			15'h000031B6 : data <= 8'b00000000 ;
			15'h000031B7 : data <= 8'b00000000 ;
			15'h000031B8 : data <= 8'b00000000 ;
			15'h000031B9 : data <= 8'b00000000 ;
			15'h000031BA : data <= 8'b00000000 ;
			15'h000031BB : data <= 8'b00000000 ;
			15'h000031BC : data <= 8'b00000000 ;
			15'h000031BD : data <= 8'b00000000 ;
			15'h000031BE : data <= 8'b00000000 ;
			15'h000031BF : data <= 8'b00000000 ;
			15'h000031C0 : data <= 8'b00000000 ;
			15'h000031C1 : data <= 8'b00000000 ;
			15'h000031C2 : data <= 8'b00000000 ;
			15'h000031C3 : data <= 8'b00000000 ;
			15'h000031C4 : data <= 8'b00000000 ;
			15'h000031C5 : data <= 8'b00000000 ;
			15'h000031C6 : data <= 8'b00000000 ;
			15'h000031C7 : data <= 8'b00000000 ;
			15'h000031C8 : data <= 8'b00000000 ;
			15'h000031C9 : data <= 8'b00000000 ;
			15'h000031CA : data <= 8'b00000000 ;
			15'h000031CB : data <= 8'b00000000 ;
			15'h000031CC : data <= 8'b00000000 ;
			15'h000031CD : data <= 8'b00000000 ;
			15'h000031CE : data <= 8'b00000000 ;
			15'h000031CF : data <= 8'b00000000 ;
			15'h000031D0 : data <= 8'b00000000 ;
			15'h000031D1 : data <= 8'b00000000 ;
			15'h000031D2 : data <= 8'b00000000 ;
			15'h000031D3 : data <= 8'b00000000 ;
			15'h000031D4 : data <= 8'b00000000 ;
			15'h000031D5 : data <= 8'b00000000 ;
			15'h000031D6 : data <= 8'b00000000 ;
			15'h000031D7 : data <= 8'b00000000 ;
			15'h000031D8 : data <= 8'b00000000 ;
			15'h000031D9 : data <= 8'b00000000 ;
			15'h000031DA : data <= 8'b00000000 ;
			15'h000031DB : data <= 8'b00000000 ;
			15'h000031DC : data <= 8'b00000000 ;
			15'h000031DD : data <= 8'b00000000 ;
			15'h000031DE : data <= 8'b00000000 ;
			15'h000031DF : data <= 8'b00000000 ;
			15'h000031E0 : data <= 8'b00000000 ;
			15'h000031E1 : data <= 8'b00000000 ;
			15'h000031E2 : data <= 8'b00000000 ;
			15'h000031E3 : data <= 8'b00000000 ;
			15'h000031E4 : data <= 8'b00000000 ;
			15'h000031E5 : data <= 8'b00000000 ;
			15'h000031E6 : data <= 8'b00000000 ;
			15'h000031E7 : data <= 8'b00000000 ;
			15'h000031E8 : data <= 8'b00000000 ;
			15'h000031E9 : data <= 8'b00000000 ;
			15'h000031EA : data <= 8'b00000000 ;
			15'h000031EB : data <= 8'b00000000 ;
			15'h000031EC : data <= 8'b00000000 ;
			15'h000031ED : data <= 8'b00000000 ;
			15'h000031EE : data <= 8'b00000000 ;
			15'h000031EF : data <= 8'b00000000 ;
			15'h000031F0 : data <= 8'b00000000 ;
			15'h000031F1 : data <= 8'b00000000 ;
			15'h000031F2 : data <= 8'b00000000 ;
			15'h000031F3 : data <= 8'b00000000 ;
			15'h000031F4 : data <= 8'b00000000 ;
			15'h000031F5 : data <= 8'b00000000 ;
			15'h000031F6 : data <= 8'b00000000 ;
			15'h000031F7 : data <= 8'b00000000 ;
			15'h000031F8 : data <= 8'b00000000 ;
			15'h000031F9 : data <= 8'b00000000 ;
			15'h000031FA : data <= 8'b00000000 ;
			15'h000031FB : data <= 8'b00000000 ;
			15'h000031FC : data <= 8'b00000000 ;
			15'h000031FD : data <= 8'b00000000 ;
			15'h000031FE : data <= 8'b00000000 ;
			15'h000031FF : data <= 8'b00000000 ;
			15'h00003200 : data <= 8'b00000000 ;
			15'h00003201 : data <= 8'b00000000 ;
			15'h00003202 : data <= 8'b00000000 ;
			15'h00003203 : data <= 8'b00000000 ;
			15'h00003204 : data <= 8'b00000000 ;
			15'h00003205 : data <= 8'b00000000 ;
			15'h00003206 : data <= 8'b00000000 ;
			15'h00003207 : data <= 8'b00000000 ;
			15'h00003208 : data <= 8'b00000000 ;
			15'h00003209 : data <= 8'b00000000 ;
			15'h0000320A : data <= 8'b00000000 ;
			15'h0000320B : data <= 8'b00000000 ;
			15'h0000320C : data <= 8'b00000000 ;
			15'h0000320D : data <= 8'b00000000 ;
			15'h0000320E : data <= 8'b00000000 ;
			15'h0000320F : data <= 8'b00000000 ;
			15'h00003210 : data <= 8'b00000000 ;
			15'h00003211 : data <= 8'b00000000 ;
			15'h00003212 : data <= 8'b00000000 ;
			15'h00003213 : data <= 8'b00000000 ;
			15'h00003214 : data <= 8'b00000000 ;
			15'h00003215 : data <= 8'b00000000 ;
			15'h00003216 : data <= 8'b00000000 ;
			15'h00003217 : data <= 8'b00000000 ;
			15'h00003218 : data <= 8'b00000000 ;
			15'h00003219 : data <= 8'b00000000 ;
			15'h0000321A : data <= 8'b00000000 ;
			15'h0000321B : data <= 8'b00000000 ;
			15'h0000321C : data <= 8'b00000000 ;
			15'h0000321D : data <= 8'b00000000 ;
			15'h0000321E : data <= 8'b00000000 ;
			15'h0000321F : data <= 8'b00000000 ;
			15'h00003220 : data <= 8'b00000000 ;
			15'h00003221 : data <= 8'b00000000 ;
			15'h00003222 : data <= 8'b00000000 ;
			15'h00003223 : data <= 8'b00000000 ;
			15'h00003224 : data <= 8'b00000000 ;
			15'h00003225 : data <= 8'b00000000 ;
			15'h00003226 : data <= 8'b00000000 ;
			15'h00003227 : data <= 8'b00000000 ;
			15'h00003228 : data <= 8'b00000000 ;
			15'h00003229 : data <= 8'b00000000 ;
			15'h0000322A : data <= 8'b00000000 ;
			15'h0000322B : data <= 8'b00000000 ;
			15'h0000322C : data <= 8'b00000000 ;
			15'h0000322D : data <= 8'b00000000 ;
			15'h0000322E : data <= 8'b00000000 ;
			15'h0000322F : data <= 8'b00000000 ;
			15'h00003230 : data <= 8'b00000000 ;
			15'h00003231 : data <= 8'b00000000 ;
			15'h00003232 : data <= 8'b00000000 ;
			15'h00003233 : data <= 8'b00000000 ;
			15'h00003234 : data <= 8'b00000000 ;
			15'h00003235 : data <= 8'b00000000 ;
			15'h00003236 : data <= 8'b00000000 ;
			15'h00003237 : data <= 8'b00000000 ;
			15'h00003238 : data <= 8'b00000000 ;
			15'h00003239 : data <= 8'b00000000 ;
			15'h0000323A : data <= 8'b00000000 ;
			15'h0000323B : data <= 8'b00000000 ;
			15'h0000323C : data <= 8'b00000000 ;
			15'h0000323D : data <= 8'b00000000 ;
			15'h0000323E : data <= 8'b00000000 ;
			15'h0000323F : data <= 8'b00000000 ;
			15'h00003240 : data <= 8'b00000000 ;
			15'h00003241 : data <= 8'b00000000 ;
			15'h00003242 : data <= 8'b00000000 ;
			15'h00003243 : data <= 8'b00000000 ;
			15'h00003244 : data <= 8'b00000000 ;
			15'h00003245 : data <= 8'b00000000 ;
			15'h00003246 : data <= 8'b00000000 ;
			15'h00003247 : data <= 8'b00000000 ;
			15'h00003248 : data <= 8'b00000000 ;
			15'h00003249 : data <= 8'b00000000 ;
			15'h0000324A : data <= 8'b00000000 ;
			15'h0000324B : data <= 8'b00000000 ;
			15'h0000324C : data <= 8'b00000000 ;
			15'h0000324D : data <= 8'b00000000 ;
			15'h0000324E : data <= 8'b00000000 ;
			15'h0000324F : data <= 8'b00000000 ;
			15'h00003250 : data <= 8'b00000000 ;
			15'h00003251 : data <= 8'b00000000 ;
			15'h00003252 : data <= 8'b00000000 ;
			15'h00003253 : data <= 8'b00000000 ;
			15'h00003254 : data <= 8'b00000000 ;
			15'h00003255 : data <= 8'b00000000 ;
			15'h00003256 : data <= 8'b00000000 ;
			15'h00003257 : data <= 8'b00000000 ;
			15'h00003258 : data <= 8'b00000000 ;
			15'h00003259 : data <= 8'b00000000 ;
			15'h0000325A : data <= 8'b00000000 ;
			15'h0000325B : data <= 8'b00000000 ;
			15'h0000325C : data <= 8'b00000000 ;
			15'h0000325D : data <= 8'b00000000 ;
			15'h0000325E : data <= 8'b00000000 ;
			15'h0000325F : data <= 8'b00000000 ;
			15'h00003260 : data <= 8'b00000000 ;
			15'h00003261 : data <= 8'b00000000 ;
			15'h00003262 : data <= 8'b00000000 ;
			15'h00003263 : data <= 8'b00000000 ;
			15'h00003264 : data <= 8'b00000000 ;
			15'h00003265 : data <= 8'b00000000 ;
			15'h00003266 : data <= 8'b00000000 ;
			15'h00003267 : data <= 8'b00000000 ;
			15'h00003268 : data <= 8'b00000000 ;
			15'h00003269 : data <= 8'b00000000 ;
			15'h0000326A : data <= 8'b00000000 ;
			15'h0000326B : data <= 8'b00000000 ;
			15'h0000326C : data <= 8'b00000000 ;
			15'h0000326D : data <= 8'b00000000 ;
			15'h0000326E : data <= 8'b00000000 ;
			15'h0000326F : data <= 8'b00000000 ;
			15'h00003270 : data <= 8'b00000000 ;
			15'h00003271 : data <= 8'b00000000 ;
			15'h00003272 : data <= 8'b00000000 ;
			15'h00003273 : data <= 8'b00000000 ;
			15'h00003274 : data <= 8'b00000000 ;
			15'h00003275 : data <= 8'b00000000 ;
			15'h00003276 : data <= 8'b00000000 ;
			15'h00003277 : data <= 8'b00000000 ;
			15'h00003278 : data <= 8'b00000000 ;
			15'h00003279 : data <= 8'b00000000 ;
			15'h0000327A : data <= 8'b00000000 ;
			15'h0000327B : data <= 8'b00000000 ;
			15'h0000327C : data <= 8'b00000000 ;
			15'h0000327D : data <= 8'b00000000 ;
			15'h0000327E : data <= 8'b00000000 ;
			15'h0000327F : data <= 8'b00000000 ;
			15'h00003280 : data <= 8'b00000000 ;
			15'h00003281 : data <= 8'b00000000 ;
			15'h00003282 : data <= 8'b00000000 ;
			15'h00003283 : data <= 8'b00000000 ;
			15'h00003284 : data <= 8'b00000000 ;
			15'h00003285 : data <= 8'b00000000 ;
			15'h00003286 : data <= 8'b00000000 ;
			15'h00003287 : data <= 8'b00000000 ;
			15'h00003288 : data <= 8'b00000000 ;
			15'h00003289 : data <= 8'b00000000 ;
			15'h0000328A : data <= 8'b00000000 ;
			15'h0000328B : data <= 8'b00000000 ;
			15'h0000328C : data <= 8'b00000000 ;
			15'h0000328D : data <= 8'b00000000 ;
			15'h0000328E : data <= 8'b00000000 ;
			15'h0000328F : data <= 8'b00000000 ;
			15'h00003290 : data <= 8'b00000000 ;
			15'h00003291 : data <= 8'b00000000 ;
			15'h00003292 : data <= 8'b00000000 ;
			15'h00003293 : data <= 8'b00000000 ;
			15'h00003294 : data <= 8'b00000000 ;
			15'h00003295 : data <= 8'b00000000 ;
			15'h00003296 : data <= 8'b00000000 ;
			15'h00003297 : data <= 8'b00000000 ;
			15'h00003298 : data <= 8'b00000000 ;
			15'h00003299 : data <= 8'b00000000 ;
			15'h0000329A : data <= 8'b00000000 ;
			15'h0000329B : data <= 8'b00000000 ;
			15'h0000329C : data <= 8'b00000000 ;
			15'h0000329D : data <= 8'b00000000 ;
			15'h0000329E : data <= 8'b00000000 ;
			15'h0000329F : data <= 8'b00000000 ;
			15'h000032A0 : data <= 8'b00000000 ;
			15'h000032A1 : data <= 8'b00000000 ;
			15'h000032A2 : data <= 8'b00000000 ;
			15'h000032A3 : data <= 8'b00000000 ;
			15'h000032A4 : data <= 8'b00000000 ;
			15'h000032A5 : data <= 8'b00000000 ;
			15'h000032A6 : data <= 8'b00000000 ;
			15'h000032A7 : data <= 8'b00000000 ;
			15'h000032A8 : data <= 8'b00000000 ;
			15'h000032A9 : data <= 8'b00000000 ;
			15'h000032AA : data <= 8'b00000000 ;
			15'h000032AB : data <= 8'b00000000 ;
			15'h000032AC : data <= 8'b00000000 ;
			15'h000032AD : data <= 8'b00000000 ;
			15'h000032AE : data <= 8'b00000000 ;
			15'h000032AF : data <= 8'b00000000 ;
			15'h000032B0 : data <= 8'b00000000 ;
			15'h000032B1 : data <= 8'b00000000 ;
			15'h000032B2 : data <= 8'b00000000 ;
			15'h000032B3 : data <= 8'b00000000 ;
			15'h000032B4 : data <= 8'b00000000 ;
			15'h000032B5 : data <= 8'b00000000 ;
			15'h000032B6 : data <= 8'b00000000 ;
			15'h000032B7 : data <= 8'b00000000 ;
			15'h000032B8 : data <= 8'b00000000 ;
			15'h000032B9 : data <= 8'b00000000 ;
			15'h000032BA : data <= 8'b00000000 ;
			15'h000032BB : data <= 8'b00000000 ;
			15'h000032BC : data <= 8'b00000000 ;
			15'h000032BD : data <= 8'b00000000 ;
			15'h000032BE : data <= 8'b00000000 ;
			15'h000032BF : data <= 8'b00000000 ;
			15'h000032C0 : data <= 8'b00000000 ;
			15'h000032C1 : data <= 8'b00000000 ;
			15'h000032C2 : data <= 8'b00000000 ;
			15'h000032C3 : data <= 8'b00000000 ;
			15'h000032C4 : data <= 8'b00000000 ;
			15'h000032C5 : data <= 8'b00000000 ;
			15'h000032C6 : data <= 8'b00000000 ;
			15'h000032C7 : data <= 8'b00000000 ;
			15'h000032C8 : data <= 8'b00000000 ;
			15'h000032C9 : data <= 8'b00000000 ;
			15'h000032CA : data <= 8'b00000000 ;
			15'h000032CB : data <= 8'b00000000 ;
			15'h000032CC : data <= 8'b00000000 ;
			15'h000032CD : data <= 8'b00000000 ;
			15'h000032CE : data <= 8'b00000000 ;
			15'h000032CF : data <= 8'b00000000 ;
			15'h000032D0 : data <= 8'b00000000 ;
			15'h000032D1 : data <= 8'b00000000 ;
			15'h000032D2 : data <= 8'b00000000 ;
			15'h000032D3 : data <= 8'b00000000 ;
			15'h000032D4 : data <= 8'b00000000 ;
			15'h000032D5 : data <= 8'b00000000 ;
			15'h000032D6 : data <= 8'b00000000 ;
			15'h000032D7 : data <= 8'b00000000 ;
			15'h000032D8 : data <= 8'b00000000 ;
			15'h000032D9 : data <= 8'b00000000 ;
			15'h000032DA : data <= 8'b00000000 ;
			15'h000032DB : data <= 8'b00000000 ;
			15'h000032DC : data <= 8'b00000000 ;
			15'h000032DD : data <= 8'b00000000 ;
			15'h000032DE : data <= 8'b00000000 ;
			15'h000032DF : data <= 8'b00000000 ;
			15'h000032E0 : data <= 8'b00000000 ;
			15'h000032E1 : data <= 8'b00000000 ;
			15'h000032E2 : data <= 8'b00000000 ;
			15'h000032E3 : data <= 8'b00000000 ;
			15'h000032E4 : data <= 8'b00000000 ;
			15'h000032E5 : data <= 8'b00000000 ;
			15'h000032E6 : data <= 8'b00000000 ;
			15'h000032E7 : data <= 8'b00000000 ;
			15'h000032E8 : data <= 8'b00000000 ;
			15'h000032E9 : data <= 8'b00000000 ;
			15'h000032EA : data <= 8'b00000000 ;
			15'h000032EB : data <= 8'b00000000 ;
			15'h000032EC : data <= 8'b00000000 ;
			15'h000032ED : data <= 8'b00000000 ;
			15'h000032EE : data <= 8'b00000000 ;
			15'h000032EF : data <= 8'b00000000 ;
			15'h000032F0 : data <= 8'b00000000 ;
			15'h000032F1 : data <= 8'b00000000 ;
			15'h000032F2 : data <= 8'b00000000 ;
			15'h000032F3 : data <= 8'b00000000 ;
			15'h000032F4 : data <= 8'b00000000 ;
			15'h000032F5 : data <= 8'b00000000 ;
			15'h000032F6 : data <= 8'b00000000 ;
			15'h000032F7 : data <= 8'b00000000 ;
			15'h000032F8 : data <= 8'b00000000 ;
			15'h000032F9 : data <= 8'b00000000 ;
			15'h000032FA : data <= 8'b00000000 ;
			15'h000032FB : data <= 8'b00000000 ;
			15'h000032FC : data <= 8'b00000000 ;
			15'h000032FD : data <= 8'b00000000 ;
			15'h000032FE : data <= 8'b00000000 ;
			15'h000032FF : data <= 8'b00000000 ;
			15'h00003300 : data <= 8'b00000000 ;
			15'h00003301 : data <= 8'b00000000 ;
			15'h00003302 : data <= 8'b00000000 ;
			15'h00003303 : data <= 8'b00000000 ;
			15'h00003304 : data <= 8'b00000000 ;
			15'h00003305 : data <= 8'b00000000 ;
			15'h00003306 : data <= 8'b00000000 ;
			15'h00003307 : data <= 8'b00000000 ;
			15'h00003308 : data <= 8'b00000000 ;
			15'h00003309 : data <= 8'b00000000 ;
			15'h0000330A : data <= 8'b00000000 ;
			15'h0000330B : data <= 8'b00000000 ;
			15'h0000330C : data <= 8'b00000000 ;
			15'h0000330D : data <= 8'b00000000 ;
			15'h0000330E : data <= 8'b00000000 ;
			15'h0000330F : data <= 8'b00000000 ;
			15'h00003310 : data <= 8'b00000000 ;
			15'h00003311 : data <= 8'b00000000 ;
			15'h00003312 : data <= 8'b00000000 ;
			15'h00003313 : data <= 8'b00000000 ;
			15'h00003314 : data <= 8'b00000000 ;
			15'h00003315 : data <= 8'b00000000 ;
			15'h00003316 : data <= 8'b00000000 ;
			15'h00003317 : data <= 8'b00000000 ;
			15'h00003318 : data <= 8'b00000000 ;
			15'h00003319 : data <= 8'b00000000 ;
			15'h0000331A : data <= 8'b00000000 ;
			15'h0000331B : data <= 8'b00000000 ;
			15'h0000331C : data <= 8'b00000000 ;
			15'h0000331D : data <= 8'b00000000 ;
			15'h0000331E : data <= 8'b00000000 ;
			15'h0000331F : data <= 8'b00000000 ;
			15'h00003320 : data <= 8'b00000000 ;
			15'h00003321 : data <= 8'b00000000 ;
			15'h00003322 : data <= 8'b00000000 ;
			15'h00003323 : data <= 8'b00000000 ;
			15'h00003324 : data <= 8'b00000000 ;
			15'h00003325 : data <= 8'b00000000 ;
			15'h00003326 : data <= 8'b00000000 ;
			15'h00003327 : data <= 8'b00000000 ;
			15'h00003328 : data <= 8'b00000000 ;
			15'h00003329 : data <= 8'b00000000 ;
			15'h0000332A : data <= 8'b00000000 ;
			15'h0000332B : data <= 8'b00000000 ;
			15'h0000332C : data <= 8'b00000000 ;
			15'h0000332D : data <= 8'b00000000 ;
			15'h0000332E : data <= 8'b00000000 ;
			15'h0000332F : data <= 8'b00000000 ;
			15'h00003330 : data <= 8'b00000000 ;
			15'h00003331 : data <= 8'b00000000 ;
			15'h00003332 : data <= 8'b00000000 ;
			15'h00003333 : data <= 8'b00000000 ;
			15'h00003334 : data <= 8'b00000000 ;
			15'h00003335 : data <= 8'b00000000 ;
			15'h00003336 : data <= 8'b00000000 ;
			15'h00003337 : data <= 8'b00000000 ;
			15'h00003338 : data <= 8'b00000000 ;
			15'h00003339 : data <= 8'b00000000 ;
			15'h0000333A : data <= 8'b00000000 ;
			15'h0000333B : data <= 8'b00000000 ;
			15'h0000333C : data <= 8'b00000000 ;
			15'h0000333D : data <= 8'b00000000 ;
			15'h0000333E : data <= 8'b00000000 ;
			15'h0000333F : data <= 8'b00000000 ;
			15'h00003340 : data <= 8'b00000000 ;
			15'h00003341 : data <= 8'b00000000 ;
			15'h00003342 : data <= 8'b00000000 ;
			15'h00003343 : data <= 8'b00000000 ;
			15'h00003344 : data <= 8'b00000000 ;
			15'h00003345 : data <= 8'b00000000 ;
			15'h00003346 : data <= 8'b00000000 ;
			15'h00003347 : data <= 8'b00000000 ;
			15'h00003348 : data <= 8'b00000000 ;
			15'h00003349 : data <= 8'b00000000 ;
			15'h0000334A : data <= 8'b00000000 ;
			15'h0000334B : data <= 8'b00000000 ;
			15'h0000334C : data <= 8'b00000000 ;
			15'h0000334D : data <= 8'b00000000 ;
			15'h0000334E : data <= 8'b00000000 ;
			15'h0000334F : data <= 8'b00000000 ;
			15'h00003350 : data <= 8'b00000000 ;
			15'h00003351 : data <= 8'b00000000 ;
			15'h00003352 : data <= 8'b00000000 ;
			15'h00003353 : data <= 8'b00000000 ;
			15'h00003354 : data <= 8'b00000000 ;
			15'h00003355 : data <= 8'b00000000 ;
			15'h00003356 : data <= 8'b00000000 ;
			15'h00003357 : data <= 8'b00000000 ;
			15'h00003358 : data <= 8'b00000000 ;
			15'h00003359 : data <= 8'b00000000 ;
			15'h0000335A : data <= 8'b00000000 ;
			15'h0000335B : data <= 8'b00000000 ;
			15'h0000335C : data <= 8'b00000000 ;
			15'h0000335D : data <= 8'b00000000 ;
			15'h0000335E : data <= 8'b00000000 ;
			15'h0000335F : data <= 8'b00000000 ;
			15'h00003360 : data <= 8'b00000000 ;
			15'h00003361 : data <= 8'b00000000 ;
			15'h00003362 : data <= 8'b00000000 ;
			15'h00003363 : data <= 8'b00000000 ;
			15'h00003364 : data <= 8'b00000000 ;
			15'h00003365 : data <= 8'b00000000 ;
			15'h00003366 : data <= 8'b00000000 ;
			15'h00003367 : data <= 8'b00000000 ;
			15'h00003368 : data <= 8'b00000000 ;
			15'h00003369 : data <= 8'b00000000 ;
			15'h0000336A : data <= 8'b00000000 ;
			15'h0000336B : data <= 8'b00000000 ;
			15'h0000336C : data <= 8'b00000000 ;
			15'h0000336D : data <= 8'b00000000 ;
			15'h0000336E : data <= 8'b00000000 ;
			15'h0000336F : data <= 8'b00000000 ;
			15'h00003370 : data <= 8'b00000000 ;
			15'h00003371 : data <= 8'b00000000 ;
			15'h00003372 : data <= 8'b00000000 ;
			15'h00003373 : data <= 8'b00000000 ;
			15'h00003374 : data <= 8'b00000000 ;
			15'h00003375 : data <= 8'b00000000 ;
			15'h00003376 : data <= 8'b00000000 ;
			15'h00003377 : data <= 8'b00000000 ;
			15'h00003378 : data <= 8'b00000000 ;
			15'h00003379 : data <= 8'b00000000 ;
			15'h0000337A : data <= 8'b00000000 ;
			15'h0000337B : data <= 8'b00000000 ;
			15'h0000337C : data <= 8'b00000000 ;
			15'h0000337D : data <= 8'b00000000 ;
			15'h0000337E : data <= 8'b00000000 ;
			15'h0000337F : data <= 8'b00000000 ;
			15'h00003380 : data <= 8'b00000000 ;
			15'h00003381 : data <= 8'b00000000 ;
			15'h00003382 : data <= 8'b00000000 ;
			15'h00003383 : data <= 8'b00000000 ;
			15'h00003384 : data <= 8'b00000000 ;
			15'h00003385 : data <= 8'b00000000 ;
			15'h00003386 : data <= 8'b00000000 ;
			15'h00003387 : data <= 8'b00000000 ;
			15'h00003388 : data <= 8'b00000000 ;
			15'h00003389 : data <= 8'b00000000 ;
			15'h0000338A : data <= 8'b00000000 ;
			15'h0000338B : data <= 8'b00000000 ;
			15'h0000338C : data <= 8'b00000000 ;
			15'h0000338D : data <= 8'b00000000 ;
			15'h0000338E : data <= 8'b00000000 ;
			15'h0000338F : data <= 8'b00000000 ;
			15'h00003390 : data <= 8'b00000000 ;
			15'h00003391 : data <= 8'b00000000 ;
			15'h00003392 : data <= 8'b00000000 ;
			15'h00003393 : data <= 8'b00000000 ;
			15'h00003394 : data <= 8'b00000000 ;
			15'h00003395 : data <= 8'b00000000 ;
			15'h00003396 : data <= 8'b00000000 ;
			15'h00003397 : data <= 8'b00000000 ;
			15'h00003398 : data <= 8'b00000000 ;
			15'h00003399 : data <= 8'b00000000 ;
			15'h0000339A : data <= 8'b00000000 ;
			15'h0000339B : data <= 8'b00000000 ;
			15'h0000339C : data <= 8'b00000000 ;
			15'h0000339D : data <= 8'b00000000 ;
			15'h0000339E : data <= 8'b00000000 ;
			15'h0000339F : data <= 8'b00000000 ;
			15'h000033A0 : data <= 8'b00000000 ;
			15'h000033A1 : data <= 8'b00000000 ;
			15'h000033A2 : data <= 8'b00000000 ;
			15'h000033A3 : data <= 8'b00000000 ;
			15'h000033A4 : data <= 8'b00000000 ;
			15'h000033A5 : data <= 8'b00000000 ;
			15'h000033A6 : data <= 8'b00000000 ;
			15'h000033A7 : data <= 8'b00000000 ;
			15'h000033A8 : data <= 8'b00000000 ;
			15'h000033A9 : data <= 8'b00000000 ;
			15'h000033AA : data <= 8'b00000000 ;
			15'h000033AB : data <= 8'b00000000 ;
			15'h000033AC : data <= 8'b00000000 ;
			15'h000033AD : data <= 8'b00000000 ;
			15'h000033AE : data <= 8'b00000000 ;
			15'h000033AF : data <= 8'b00000000 ;
			15'h000033B0 : data <= 8'b00000000 ;
			15'h000033B1 : data <= 8'b00000000 ;
			15'h000033B2 : data <= 8'b00000000 ;
			15'h000033B3 : data <= 8'b00000000 ;
			15'h000033B4 : data <= 8'b00000000 ;
			15'h000033B5 : data <= 8'b00000000 ;
			15'h000033B6 : data <= 8'b00000000 ;
			15'h000033B7 : data <= 8'b00000000 ;
			15'h000033B8 : data <= 8'b00000000 ;
			15'h000033B9 : data <= 8'b00000000 ;
			15'h000033BA : data <= 8'b00000000 ;
			15'h000033BB : data <= 8'b00000000 ;
			15'h000033BC : data <= 8'b00000000 ;
			15'h000033BD : data <= 8'b00000000 ;
			15'h000033BE : data <= 8'b00000000 ;
			15'h000033BF : data <= 8'b00000000 ;
			15'h000033C0 : data <= 8'b00000000 ;
			15'h000033C1 : data <= 8'b00000000 ;
			15'h000033C2 : data <= 8'b00000000 ;
			15'h000033C3 : data <= 8'b00000000 ;
			15'h000033C4 : data <= 8'b00000000 ;
			15'h000033C5 : data <= 8'b00000000 ;
			15'h000033C6 : data <= 8'b00000000 ;
			15'h000033C7 : data <= 8'b00000000 ;
			15'h000033C8 : data <= 8'b00000000 ;
			15'h000033C9 : data <= 8'b00000000 ;
			15'h000033CA : data <= 8'b00000000 ;
			15'h000033CB : data <= 8'b00000000 ;
			15'h000033CC : data <= 8'b00000000 ;
			15'h000033CD : data <= 8'b00000000 ;
			15'h000033CE : data <= 8'b00000000 ;
			15'h000033CF : data <= 8'b00000000 ;
			15'h000033D0 : data <= 8'b00000000 ;
			15'h000033D1 : data <= 8'b00000000 ;
			15'h000033D2 : data <= 8'b00000000 ;
			15'h000033D3 : data <= 8'b00000000 ;
			15'h000033D4 : data <= 8'b00000000 ;
			15'h000033D5 : data <= 8'b00000000 ;
			15'h000033D6 : data <= 8'b00000000 ;
			15'h000033D7 : data <= 8'b00000000 ;
			15'h000033D8 : data <= 8'b00000000 ;
			15'h000033D9 : data <= 8'b00000000 ;
			15'h000033DA : data <= 8'b00000000 ;
			15'h000033DB : data <= 8'b00000000 ;
			15'h000033DC : data <= 8'b00000000 ;
			15'h000033DD : data <= 8'b00000000 ;
			15'h000033DE : data <= 8'b00000000 ;
			15'h000033DF : data <= 8'b00000000 ;
			15'h000033E0 : data <= 8'b00000000 ;
			15'h000033E1 : data <= 8'b00000000 ;
			15'h000033E2 : data <= 8'b00000000 ;
			15'h000033E3 : data <= 8'b00000000 ;
			15'h000033E4 : data <= 8'b00000000 ;
			15'h000033E5 : data <= 8'b00000000 ;
			15'h000033E6 : data <= 8'b00000000 ;
			15'h000033E7 : data <= 8'b00000000 ;
			15'h000033E8 : data <= 8'b00000000 ;
			15'h000033E9 : data <= 8'b00000000 ;
			15'h000033EA : data <= 8'b00000000 ;
			15'h000033EB : data <= 8'b00000000 ;
			15'h000033EC : data <= 8'b00000000 ;
			15'h000033ED : data <= 8'b00000000 ;
			15'h000033EE : data <= 8'b00000000 ;
			15'h000033EF : data <= 8'b00000000 ;
			15'h000033F0 : data <= 8'b00000000 ;
			15'h000033F1 : data <= 8'b00000000 ;
			15'h000033F2 : data <= 8'b00000000 ;
			15'h000033F3 : data <= 8'b00000000 ;
			15'h000033F4 : data <= 8'b00000000 ;
			15'h000033F5 : data <= 8'b00000000 ;
			15'h000033F6 : data <= 8'b00000000 ;
			15'h000033F7 : data <= 8'b00000000 ;
			15'h000033F8 : data <= 8'b00000000 ;
			15'h000033F9 : data <= 8'b00000000 ;
			15'h000033FA : data <= 8'b00000000 ;
			15'h000033FB : data <= 8'b00000000 ;
			15'h000033FC : data <= 8'b00000000 ;
			15'h000033FD : data <= 8'b00000000 ;
			15'h000033FE : data <= 8'b00000000 ;
			15'h000033FF : data <= 8'b00000000 ;
			15'h00003400 : data <= 8'b00000000 ;
			15'h00003401 : data <= 8'b00000000 ;
			15'h00003402 : data <= 8'b00000000 ;
			15'h00003403 : data <= 8'b00000000 ;
			15'h00003404 : data <= 8'b00000000 ;
			15'h00003405 : data <= 8'b00000000 ;
			15'h00003406 : data <= 8'b00000000 ;
			15'h00003407 : data <= 8'b00000000 ;
			15'h00003408 : data <= 8'b00000000 ;
			15'h00003409 : data <= 8'b00000000 ;
			15'h0000340A : data <= 8'b00000000 ;
			15'h0000340B : data <= 8'b00000000 ;
			15'h0000340C : data <= 8'b00000000 ;
			15'h0000340D : data <= 8'b00000000 ;
			15'h0000340E : data <= 8'b00000000 ;
			15'h0000340F : data <= 8'b00000000 ;
			15'h00003410 : data <= 8'b00000000 ;
			15'h00003411 : data <= 8'b00000000 ;
			15'h00003412 : data <= 8'b00000000 ;
			15'h00003413 : data <= 8'b00000000 ;
			15'h00003414 : data <= 8'b00000000 ;
			15'h00003415 : data <= 8'b00000000 ;
			15'h00003416 : data <= 8'b00000000 ;
			15'h00003417 : data <= 8'b00000000 ;
			15'h00003418 : data <= 8'b00000000 ;
			15'h00003419 : data <= 8'b00000000 ;
			15'h0000341A : data <= 8'b00000000 ;
			15'h0000341B : data <= 8'b00000000 ;
			15'h0000341C : data <= 8'b00000000 ;
			15'h0000341D : data <= 8'b00000000 ;
			15'h0000341E : data <= 8'b00000000 ;
			15'h0000341F : data <= 8'b00000000 ;
			15'h00003420 : data <= 8'b00000000 ;
			15'h00003421 : data <= 8'b00000000 ;
			15'h00003422 : data <= 8'b00000000 ;
			15'h00003423 : data <= 8'b00000000 ;
			15'h00003424 : data <= 8'b00000000 ;
			15'h00003425 : data <= 8'b00000000 ;
			15'h00003426 : data <= 8'b00000000 ;
			15'h00003427 : data <= 8'b00000000 ;
			15'h00003428 : data <= 8'b00000000 ;
			15'h00003429 : data <= 8'b00000000 ;
			15'h0000342A : data <= 8'b00000000 ;
			15'h0000342B : data <= 8'b00000000 ;
			15'h0000342C : data <= 8'b00000000 ;
			15'h0000342D : data <= 8'b00000000 ;
			15'h0000342E : data <= 8'b00000000 ;
			15'h0000342F : data <= 8'b00000000 ;
			15'h00003430 : data <= 8'b00000000 ;
			15'h00003431 : data <= 8'b00000000 ;
			15'h00003432 : data <= 8'b00000000 ;
			15'h00003433 : data <= 8'b00000000 ;
			15'h00003434 : data <= 8'b00000000 ;
			15'h00003435 : data <= 8'b00000000 ;
			15'h00003436 : data <= 8'b00000000 ;
			15'h00003437 : data <= 8'b00000000 ;
			15'h00003438 : data <= 8'b00000000 ;
			15'h00003439 : data <= 8'b00000000 ;
			15'h0000343A : data <= 8'b00000000 ;
			15'h0000343B : data <= 8'b00000000 ;
			15'h0000343C : data <= 8'b00000000 ;
			15'h0000343D : data <= 8'b00000000 ;
			15'h0000343E : data <= 8'b00000000 ;
			15'h0000343F : data <= 8'b00000000 ;
			15'h00003440 : data <= 8'b00000000 ;
			15'h00003441 : data <= 8'b00000000 ;
			15'h00003442 : data <= 8'b00000000 ;
			15'h00003443 : data <= 8'b00000000 ;
			15'h00003444 : data <= 8'b00000000 ;
			15'h00003445 : data <= 8'b00000000 ;
			15'h00003446 : data <= 8'b00000000 ;
			15'h00003447 : data <= 8'b00000000 ;
			15'h00003448 : data <= 8'b00000000 ;
			15'h00003449 : data <= 8'b00000000 ;
			15'h0000344A : data <= 8'b00000000 ;
			15'h0000344B : data <= 8'b00000000 ;
			15'h0000344C : data <= 8'b00000000 ;
			15'h0000344D : data <= 8'b00000000 ;
			15'h0000344E : data <= 8'b00000000 ;
			15'h0000344F : data <= 8'b00000000 ;
			15'h00003450 : data <= 8'b00000000 ;
			15'h00003451 : data <= 8'b00000000 ;
			15'h00003452 : data <= 8'b00000000 ;
			15'h00003453 : data <= 8'b00000000 ;
			15'h00003454 : data <= 8'b00000000 ;
			15'h00003455 : data <= 8'b00000000 ;
			15'h00003456 : data <= 8'b00000000 ;
			15'h00003457 : data <= 8'b00000000 ;
			15'h00003458 : data <= 8'b00000000 ;
			15'h00003459 : data <= 8'b00000000 ;
			15'h0000345A : data <= 8'b00000000 ;
			15'h0000345B : data <= 8'b00000000 ;
			15'h0000345C : data <= 8'b00000000 ;
			15'h0000345D : data <= 8'b00000000 ;
			15'h0000345E : data <= 8'b00000000 ;
			15'h0000345F : data <= 8'b00000000 ;
			15'h00003460 : data <= 8'b00000000 ;
			15'h00003461 : data <= 8'b00000000 ;
			15'h00003462 : data <= 8'b00000000 ;
			15'h00003463 : data <= 8'b00000000 ;
			15'h00003464 : data <= 8'b00000000 ;
			15'h00003465 : data <= 8'b00000000 ;
			15'h00003466 : data <= 8'b00000000 ;
			15'h00003467 : data <= 8'b00000000 ;
			15'h00003468 : data <= 8'b00000000 ;
			15'h00003469 : data <= 8'b00000000 ;
			15'h0000346A : data <= 8'b00000000 ;
			15'h0000346B : data <= 8'b00000000 ;
			15'h0000346C : data <= 8'b00000000 ;
			15'h0000346D : data <= 8'b00000000 ;
			15'h0000346E : data <= 8'b00000000 ;
			15'h0000346F : data <= 8'b00000000 ;
			15'h00003470 : data <= 8'b00000000 ;
			15'h00003471 : data <= 8'b00000000 ;
			15'h00003472 : data <= 8'b00000000 ;
			15'h00003473 : data <= 8'b00000000 ;
			15'h00003474 : data <= 8'b00000000 ;
			15'h00003475 : data <= 8'b00000000 ;
			15'h00003476 : data <= 8'b00000000 ;
			15'h00003477 : data <= 8'b00000000 ;
			15'h00003478 : data <= 8'b00000000 ;
			15'h00003479 : data <= 8'b00000000 ;
			15'h0000347A : data <= 8'b00000000 ;
			15'h0000347B : data <= 8'b00000000 ;
			15'h0000347C : data <= 8'b00000000 ;
			15'h0000347D : data <= 8'b00000000 ;
			15'h0000347E : data <= 8'b00000000 ;
			15'h0000347F : data <= 8'b00000000 ;
			15'h00003480 : data <= 8'b00000000 ;
			15'h00003481 : data <= 8'b00000000 ;
			15'h00003482 : data <= 8'b00000000 ;
			15'h00003483 : data <= 8'b00000000 ;
			15'h00003484 : data <= 8'b00000000 ;
			15'h00003485 : data <= 8'b00000000 ;
			15'h00003486 : data <= 8'b00000000 ;
			15'h00003487 : data <= 8'b00000000 ;
			15'h00003488 : data <= 8'b00000000 ;
			15'h00003489 : data <= 8'b00000000 ;
			15'h0000348A : data <= 8'b00000000 ;
			15'h0000348B : data <= 8'b00000000 ;
			15'h0000348C : data <= 8'b00000000 ;
			15'h0000348D : data <= 8'b00000000 ;
			15'h0000348E : data <= 8'b00000000 ;
			15'h0000348F : data <= 8'b00000000 ;
			15'h00003490 : data <= 8'b00000000 ;
			15'h00003491 : data <= 8'b00000000 ;
			15'h00003492 : data <= 8'b00000000 ;
			15'h00003493 : data <= 8'b00000000 ;
			15'h00003494 : data <= 8'b00000000 ;
			15'h00003495 : data <= 8'b00000000 ;
			15'h00003496 : data <= 8'b00000000 ;
			15'h00003497 : data <= 8'b00000000 ;
			15'h00003498 : data <= 8'b00000000 ;
			15'h00003499 : data <= 8'b00000000 ;
			15'h0000349A : data <= 8'b00000000 ;
			15'h0000349B : data <= 8'b00000000 ;
			15'h0000349C : data <= 8'b00000000 ;
			15'h0000349D : data <= 8'b00000000 ;
			15'h0000349E : data <= 8'b00000000 ;
			15'h0000349F : data <= 8'b00000000 ;
			15'h000034A0 : data <= 8'b00000000 ;
			15'h000034A1 : data <= 8'b00000000 ;
			15'h000034A2 : data <= 8'b00000000 ;
			15'h000034A3 : data <= 8'b00000000 ;
			15'h000034A4 : data <= 8'b00000000 ;
			15'h000034A5 : data <= 8'b00000000 ;
			15'h000034A6 : data <= 8'b00000000 ;
			15'h000034A7 : data <= 8'b00000000 ;
			15'h000034A8 : data <= 8'b00000000 ;
			15'h000034A9 : data <= 8'b00000000 ;
			15'h000034AA : data <= 8'b00000000 ;
			15'h000034AB : data <= 8'b00000000 ;
			15'h000034AC : data <= 8'b00000000 ;
			15'h000034AD : data <= 8'b00000000 ;
			15'h000034AE : data <= 8'b00000000 ;
			15'h000034AF : data <= 8'b00000000 ;
			15'h000034B0 : data <= 8'b00000000 ;
			15'h000034B1 : data <= 8'b00000000 ;
			15'h000034B2 : data <= 8'b00000000 ;
			15'h000034B3 : data <= 8'b00000000 ;
			15'h000034B4 : data <= 8'b00000000 ;
			15'h000034B5 : data <= 8'b00000000 ;
			15'h000034B6 : data <= 8'b00000000 ;
			15'h000034B7 : data <= 8'b00000000 ;
			15'h000034B8 : data <= 8'b00000000 ;
			15'h000034B9 : data <= 8'b00000000 ;
			15'h000034BA : data <= 8'b00000000 ;
			15'h000034BB : data <= 8'b00000000 ;
			15'h000034BC : data <= 8'b00000000 ;
			15'h000034BD : data <= 8'b00000000 ;
			15'h000034BE : data <= 8'b00000000 ;
			15'h000034BF : data <= 8'b00000000 ;
			15'h000034C0 : data <= 8'b00000000 ;
			15'h000034C1 : data <= 8'b00000000 ;
			15'h000034C2 : data <= 8'b00000000 ;
			15'h000034C3 : data <= 8'b00000000 ;
			15'h000034C4 : data <= 8'b00000000 ;
			15'h000034C5 : data <= 8'b00000000 ;
			15'h000034C6 : data <= 8'b00000000 ;
			15'h000034C7 : data <= 8'b00000000 ;
			15'h000034C8 : data <= 8'b00000000 ;
			15'h000034C9 : data <= 8'b00000000 ;
			15'h000034CA : data <= 8'b00000000 ;
			15'h000034CB : data <= 8'b00000000 ;
			15'h000034CC : data <= 8'b00000000 ;
			15'h000034CD : data <= 8'b00000000 ;
			15'h000034CE : data <= 8'b00000000 ;
			15'h000034CF : data <= 8'b00000000 ;
			15'h000034D0 : data <= 8'b00000000 ;
			15'h000034D1 : data <= 8'b00000000 ;
			15'h000034D2 : data <= 8'b00000000 ;
			15'h000034D3 : data <= 8'b00000000 ;
			15'h000034D4 : data <= 8'b00000000 ;
			15'h000034D5 : data <= 8'b00000000 ;
			15'h000034D6 : data <= 8'b00000000 ;
			15'h000034D7 : data <= 8'b00000000 ;
			15'h000034D8 : data <= 8'b00000000 ;
			15'h000034D9 : data <= 8'b00000000 ;
			15'h000034DA : data <= 8'b00000000 ;
			15'h000034DB : data <= 8'b00000000 ;
			15'h000034DC : data <= 8'b00000000 ;
			15'h000034DD : data <= 8'b00000000 ;
			15'h000034DE : data <= 8'b00000000 ;
			15'h000034DF : data <= 8'b00000000 ;
			15'h000034E0 : data <= 8'b00000000 ;
			15'h000034E1 : data <= 8'b00000000 ;
			15'h000034E2 : data <= 8'b00000000 ;
			15'h000034E3 : data <= 8'b00000000 ;
			15'h000034E4 : data <= 8'b00000000 ;
			15'h000034E5 : data <= 8'b00000000 ;
			15'h000034E6 : data <= 8'b00000000 ;
			15'h000034E7 : data <= 8'b00000000 ;
			15'h000034E8 : data <= 8'b00000000 ;
			15'h000034E9 : data <= 8'b00000000 ;
			15'h000034EA : data <= 8'b00000000 ;
			15'h000034EB : data <= 8'b00000000 ;
			15'h000034EC : data <= 8'b00000000 ;
			15'h000034ED : data <= 8'b00000000 ;
			15'h000034EE : data <= 8'b00000000 ;
			15'h000034EF : data <= 8'b00000000 ;
			15'h000034F0 : data <= 8'b00000000 ;
			15'h000034F1 : data <= 8'b00000000 ;
			15'h000034F2 : data <= 8'b00000000 ;
			15'h000034F3 : data <= 8'b00000000 ;
			15'h000034F4 : data <= 8'b00000000 ;
			15'h000034F5 : data <= 8'b00000000 ;
			15'h000034F6 : data <= 8'b00000000 ;
			15'h000034F7 : data <= 8'b00000000 ;
			15'h000034F8 : data <= 8'b00000000 ;
			15'h000034F9 : data <= 8'b00000000 ;
			15'h000034FA : data <= 8'b00000000 ;
			15'h000034FB : data <= 8'b00000000 ;
			15'h000034FC : data <= 8'b00000000 ;
			15'h000034FD : data <= 8'b00000000 ;
			15'h000034FE : data <= 8'b00000000 ;
			15'h000034FF : data <= 8'b00000000 ;
			15'h00003500 : data <= 8'b00000000 ;
			15'h00003501 : data <= 8'b00000000 ;
			15'h00003502 : data <= 8'b00000000 ;
			15'h00003503 : data <= 8'b00000000 ;
			15'h00003504 : data <= 8'b00000000 ;
			15'h00003505 : data <= 8'b00000000 ;
			15'h00003506 : data <= 8'b00000000 ;
			15'h00003507 : data <= 8'b00000000 ;
			15'h00003508 : data <= 8'b00000000 ;
			15'h00003509 : data <= 8'b00000000 ;
			15'h0000350A : data <= 8'b00000000 ;
			15'h0000350B : data <= 8'b00000000 ;
			15'h0000350C : data <= 8'b00000000 ;
			15'h0000350D : data <= 8'b00000000 ;
			15'h0000350E : data <= 8'b00000000 ;
			15'h0000350F : data <= 8'b00000000 ;
			15'h00003510 : data <= 8'b00000000 ;
			15'h00003511 : data <= 8'b00000000 ;
			15'h00003512 : data <= 8'b00000000 ;
			15'h00003513 : data <= 8'b00000000 ;
			15'h00003514 : data <= 8'b00000000 ;
			15'h00003515 : data <= 8'b00000000 ;
			15'h00003516 : data <= 8'b00000000 ;
			15'h00003517 : data <= 8'b00000000 ;
			15'h00003518 : data <= 8'b00000000 ;
			15'h00003519 : data <= 8'b00000000 ;
			15'h0000351A : data <= 8'b00000000 ;
			15'h0000351B : data <= 8'b00000000 ;
			15'h0000351C : data <= 8'b00000000 ;
			15'h0000351D : data <= 8'b00000000 ;
			15'h0000351E : data <= 8'b00000000 ;
			15'h0000351F : data <= 8'b00000000 ;
			15'h00003520 : data <= 8'b00000000 ;
			15'h00003521 : data <= 8'b00000000 ;
			15'h00003522 : data <= 8'b00000000 ;
			15'h00003523 : data <= 8'b00000000 ;
			15'h00003524 : data <= 8'b00000000 ;
			15'h00003525 : data <= 8'b00000000 ;
			15'h00003526 : data <= 8'b00000000 ;
			15'h00003527 : data <= 8'b00000000 ;
			15'h00003528 : data <= 8'b00000000 ;
			15'h00003529 : data <= 8'b00000000 ;
			15'h0000352A : data <= 8'b00000000 ;
			15'h0000352B : data <= 8'b00000000 ;
			15'h0000352C : data <= 8'b00000000 ;
			15'h0000352D : data <= 8'b00000000 ;
			15'h0000352E : data <= 8'b00000000 ;
			15'h0000352F : data <= 8'b00000000 ;
			15'h00003530 : data <= 8'b00000000 ;
			15'h00003531 : data <= 8'b00000000 ;
			15'h00003532 : data <= 8'b00000000 ;
			15'h00003533 : data <= 8'b00000000 ;
			15'h00003534 : data <= 8'b00000000 ;
			15'h00003535 : data <= 8'b00000000 ;
			15'h00003536 : data <= 8'b00000000 ;
			15'h00003537 : data <= 8'b00000000 ;
			15'h00003538 : data <= 8'b00000000 ;
			15'h00003539 : data <= 8'b00000000 ;
			15'h0000353A : data <= 8'b00000000 ;
			15'h0000353B : data <= 8'b00000000 ;
			15'h0000353C : data <= 8'b00000000 ;
			15'h0000353D : data <= 8'b00000000 ;
			15'h0000353E : data <= 8'b00000000 ;
			15'h0000353F : data <= 8'b00000000 ;
			15'h00003540 : data <= 8'b00000000 ;
			15'h00003541 : data <= 8'b00000000 ;
			15'h00003542 : data <= 8'b00000000 ;
			15'h00003543 : data <= 8'b00000000 ;
			15'h00003544 : data <= 8'b00000000 ;
			15'h00003545 : data <= 8'b00000000 ;
			15'h00003546 : data <= 8'b00000000 ;
			15'h00003547 : data <= 8'b00000000 ;
			15'h00003548 : data <= 8'b00000000 ;
			15'h00003549 : data <= 8'b00000000 ;
			15'h0000354A : data <= 8'b00000000 ;
			15'h0000354B : data <= 8'b00000000 ;
			15'h0000354C : data <= 8'b00000000 ;
			15'h0000354D : data <= 8'b00000000 ;
			15'h0000354E : data <= 8'b00000000 ;
			15'h0000354F : data <= 8'b00000000 ;
			15'h00003550 : data <= 8'b00000000 ;
			15'h00003551 : data <= 8'b00000000 ;
			15'h00003552 : data <= 8'b00000000 ;
			15'h00003553 : data <= 8'b00000000 ;
			15'h00003554 : data <= 8'b00000000 ;
			15'h00003555 : data <= 8'b00000000 ;
			15'h00003556 : data <= 8'b00000000 ;
			15'h00003557 : data <= 8'b00000000 ;
			15'h00003558 : data <= 8'b00000000 ;
			15'h00003559 : data <= 8'b00000000 ;
			15'h0000355A : data <= 8'b00000000 ;
			15'h0000355B : data <= 8'b00000000 ;
			15'h0000355C : data <= 8'b00000000 ;
			15'h0000355D : data <= 8'b00000000 ;
			15'h0000355E : data <= 8'b00000000 ;
			15'h0000355F : data <= 8'b00000000 ;
			15'h00003560 : data <= 8'b00000000 ;
			15'h00003561 : data <= 8'b00000000 ;
			15'h00003562 : data <= 8'b00000000 ;
			15'h00003563 : data <= 8'b00000000 ;
			15'h00003564 : data <= 8'b00000000 ;
			15'h00003565 : data <= 8'b00000000 ;
			15'h00003566 : data <= 8'b00000000 ;
			15'h00003567 : data <= 8'b00000000 ;
			15'h00003568 : data <= 8'b00000000 ;
			15'h00003569 : data <= 8'b00000000 ;
			15'h0000356A : data <= 8'b00000000 ;
			15'h0000356B : data <= 8'b00000000 ;
			15'h0000356C : data <= 8'b00000000 ;
			15'h0000356D : data <= 8'b00000000 ;
			15'h0000356E : data <= 8'b00000000 ;
			15'h0000356F : data <= 8'b00000000 ;
			15'h00003570 : data <= 8'b00000000 ;
			15'h00003571 : data <= 8'b00000000 ;
			15'h00003572 : data <= 8'b00000000 ;
			15'h00003573 : data <= 8'b00000000 ;
			15'h00003574 : data <= 8'b00000000 ;
			15'h00003575 : data <= 8'b00000000 ;
			15'h00003576 : data <= 8'b00000000 ;
			15'h00003577 : data <= 8'b00000000 ;
			15'h00003578 : data <= 8'b00000000 ;
			15'h00003579 : data <= 8'b00000000 ;
			15'h0000357A : data <= 8'b00000000 ;
			15'h0000357B : data <= 8'b00000000 ;
			15'h0000357C : data <= 8'b00000000 ;
			15'h0000357D : data <= 8'b00000000 ;
			15'h0000357E : data <= 8'b00000000 ;
			15'h0000357F : data <= 8'b00000000 ;
			15'h00003580 : data <= 8'b00000000 ;
			15'h00003581 : data <= 8'b00000000 ;
			15'h00003582 : data <= 8'b00000000 ;
			15'h00003583 : data <= 8'b00000000 ;
			15'h00003584 : data <= 8'b00000000 ;
			15'h00003585 : data <= 8'b00000000 ;
			15'h00003586 : data <= 8'b00000000 ;
			15'h00003587 : data <= 8'b00000000 ;
			15'h00003588 : data <= 8'b00000000 ;
			15'h00003589 : data <= 8'b00000000 ;
			15'h0000358A : data <= 8'b00000000 ;
			15'h0000358B : data <= 8'b00000000 ;
			15'h0000358C : data <= 8'b00000000 ;
			15'h0000358D : data <= 8'b00000000 ;
			15'h0000358E : data <= 8'b00000000 ;
			15'h0000358F : data <= 8'b00000000 ;
			15'h00003590 : data <= 8'b00000000 ;
			15'h00003591 : data <= 8'b00000000 ;
			15'h00003592 : data <= 8'b00000000 ;
			15'h00003593 : data <= 8'b00000000 ;
			15'h00003594 : data <= 8'b00000000 ;
			15'h00003595 : data <= 8'b00000000 ;
			15'h00003596 : data <= 8'b00000000 ;
			15'h00003597 : data <= 8'b00000000 ;
			15'h00003598 : data <= 8'b00000000 ;
			15'h00003599 : data <= 8'b00000000 ;
			15'h0000359A : data <= 8'b00000000 ;
			15'h0000359B : data <= 8'b00000000 ;
			15'h0000359C : data <= 8'b00000000 ;
			15'h0000359D : data <= 8'b00000000 ;
			15'h0000359E : data <= 8'b00000000 ;
			15'h0000359F : data <= 8'b00000000 ;
			15'h000035A0 : data <= 8'b00000000 ;
			15'h000035A1 : data <= 8'b00000000 ;
			15'h000035A2 : data <= 8'b00000000 ;
			15'h000035A3 : data <= 8'b00000000 ;
			15'h000035A4 : data <= 8'b00000000 ;
			15'h000035A5 : data <= 8'b00000000 ;
			15'h000035A6 : data <= 8'b00000000 ;
			15'h000035A7 : data <= 8'b00000000 ;
			15'h000035A8 : data <= 8'b00000000 ;
			15'h000035A9 : data <= 8'b00000000 ;
			15'h000035AA : data <= 8'b00000000 ;
			15'h000035AB : data <= 8'b00000000 ;
			15'h000035AC : data <= 8'b00000000 ;
			15'h000035AD : data <= 8'b00000000 ;
			15'h000035AE : data <= 8'b00000000 ;
			15'h000035AF : data <= 8'b00000000 ;
			15'h000035B0 : data <= 8'b00000000 ;
			15'h000035B1 : data <= 8'b00000000 ;
			15'h000035B2 : data <= 8'b00000000 ;
			15'h000035B3 : data <= 8'b00000000 ;
			15'h000035B4 : data <= 8'b00000000 ;
			15'h000035B5 : data <= 8'b00000000 ;
			15'h000035B6 : data <= 8'b00000000 ;
			15'h000035B7 : data <= 8'b00000000 ;
			15'h000035B8 : data <= 8'b00000000 ;
			15'h000035B9 : data <= 8'b00000000 ;
			15'h000035BA : data <= 8'b00000000 ;
			15'h000035BB : data <= 8'b00000000 ;
			15'h000035BC : data <= 8'b00000000 ;
			15'h000035BD : data <= 8'b00000000 ;
			15'h000035BE : data <= 8'b00000000 ;
			15'h000035BF : data <= 8'b00000000 ;
			15'h000035C0 : data <= 8'b00000000 ;
			15'h000035C1 : data <= 8'b00000000 ;
			15'h000035C2 : data <= 8'b00000000 ;
			15'h000035C3 : data <= 8'b00000000 ;
			15'h000035C4 : data <= 8'b00000000 ;
			15'h000035C5 : data <= 8'b00000000 ;
			15'h000035C6 : data <= 8'b00000000 ;
			15'h000035C7 : data <= 8'b00000000 ;
			15'h000035C8 : data <= 8'b00000000 ;
			15'h000035C9 : data <= 8'b00000000 ;
			15'h000035CA : data <= 8'b00000000 ;
			15'h000035CB : data <= 8'b00000000 ;
			15'h000035CC : data <= 8'b00000000 ;
			15'h000035CD : data <= 8'b00000000 ;
			15'h000035CE : data <= 8'b00000000 ;
			15'h000035CF : data <= 8'b00000000 ;
			15'h000035D0 : data <= 8'b00000000 ;
			15'h000035D1 : data <= 8'b00000000 ;
			15'h000035D2 : data <= 8'b00000000 ;
			15'h000035D3 : data <= 8'b00000000 ;
			15'h000035D4 : data <= 8'b00000000 ;
			15'h000035D5 : data <= 8'b00000000 ;
			15'h000035D6 : data <= 8'b00000000 ;
			15'h000035D7 : data <= 8'b00000000 ;
			15'h000035D8 : data <= 8'b00000000 ;
			15'h000035D9 : data <= 8'b00000000 ;
			15'h000035DA : data <= 8'b00000000 ;
			15'h000035DB : data <= 8'b00000000 ;
			15'h000035DC : data <= 8'b00000000 ;
			15'h000035DD : data <= 8'b00000000 ;
			15'h000035DE : data <= 8'b00000000 ;
			15'h000035DF : data <= 8'b00000000 ;
			15'h000035E0 : data <= 8'b00000000 ;
			15'h000035E1 : data <= 8'b00000000 ;
			15'h000035E2 : data <= 8'b00000000 ;
			15'h000035E3 : data <= 8'b00000000 ;
			15'h000035E4 : data <= 8'b00000000 ;
			15'h000035E5 : data <= 8'b00000000 ;
			15'h000035E6 : data <= 8'b00000000 ;
			15'h000035E7 : data <= 8'b00000000 ;
			15'h000035E8 : data <= 8'b00000000 ;
			15'h000035E9 : data <= 8'b00000000 ;
			15'h000035EA : data <= 8'b00000000 ;
			15'h000035EB : data <= 8'b00000000 ;
			15'h000035EC : data <= 8'b00000000 ;
			15'h000035ED : data <= 8'b00000000 ;
			15'h000035EE : data <= 8'b00000000 ;
			15'h000035EF : data <= 8'b00000000 ;
			15'h000035F0 : data <= 8'b00000000 ;
			15'h000035F1 : data <= 8'b00000000 ;
			15'h000035F2 : data <= 8'b00000000 ;
			15'h000035F3 : data <= 8'b00000000 ;
			15'h000035F4 : data <= 8'b00000000 ;
			15'h000035F5 : data <= 8'b00000000 ;
			15'h000035F6 : data <= 8'b00000000 ;
			15'h000035F7 : data <= 8'b00000000 ;
			15'h000035F8 : data <= 8'b00000000 ;
			15'h000035F9 : data <= 8'b00000000 ;
			15'h000035FA : data <= 8'b00000000 ;
			15'h000035FB : data <= 8'b00000000 ;
			15'h000035FC : data <= 8'b00000000 ;
			15'h000035FD : data <= 8'b00000000 ;
			15'h000035FE : data <= 8'b00000000 ;
			15'h000035FF : data <= 8'b00000000 ;
			15'h00003600 : data <= 8'b00000000 ;
			15'h00003601 : data <= 8'b00000000 ;
			15'h00003602 : data <= 8'b00000000 ;
			15'h00003603 : data <= 8'b00000000 ;
			15'h00003604 : data <= 8'b00000000 ;
			15'h00003605 : data <= 8'b00000000 ;
			15'h00003606 : data <= 8'b00000000 ;
			15'h00003607 : data <= 8'b00000000 ;
			15'h00003608 : data <= 8'b00000000 ;
			15'h00003609 : data <= 8'b00000000 ;
			15'h0000360A : data <= 8'b00000000 ;
			15'h0000360B : data <= 8'b00000000 ;
			15'h0000360C : data <= 8'b00000000 ;
			15'h0000360D : data <= 8'b00000000 ;
			15'h0000360E : data <= 8'b00000000 ;
			15'h0000360F : data <= 8'b00000000 ;
			15'h00003610 : data <= 8'b00000000 ;
			15'h00003611 : data <= 8'b00000000 ;
			15'h00003612 : data <= 8'b00000000 ;
			15'h00003613 : data <= 8'b00000000 ;
			15'h00003614 : data <= 8'b00000000 ;
			15'h00003615 : data <= 8'b00000000 ;
			15'h00003616 : data <= 8'b00000000 ;
			15'h00003617 : data <= 8'b00000000 ;
			15'h00003618 : data <= 8'b00000000 ;
			15'h00003619 : data <= 8'b00000000 ;
			15'h0000361A : data <= 8'b00000000 ;
			15'h0000361B : data <= 8'b00000000 ;
			15'h0000361C : data <= 8'b00000000 ;
			15'h0000361D : data <= 8'b00000000 ;
			15'h0000361E : data <= 8'b00000000 ;
			15'h0000361F : data <= 8'b00000000 ;
			15'h00003620 : data <= 8'b00000000 ;
			15'h00003621 : data <= 8'b00000000 ;
			15'h00003622 : data <= 8'b00000000 ;
			15'h00003623 : data <= 8'b00000000 ;
			15'h00003624 : data <= 8'b00000000 ;
			15'h00003625 : data <= 8'b00000000 ;
			15'h00003626 : data <= 8'b00000000 ;
			15'h00003627 : data <= 8'b00000000 ;
			15'h00003628 : data <= 8'b00000000 ;
			15'h00003629 : data <= 8'b00000000 ;
			15'h0000362A : data <= 8'b00000000 ;
			15'h0000362B : data <= 8'b00000000 ;
			15'h0000362C : data <= 8'b00000000 ;
			15'h0000362D : data <= 8'b00000000 ;
			15'h0000362E : data <= 8'b00000000 ;
			15'h0000362F : data <= 8'b00000000 ;
			15'h00003630 : data <= 8'b00000000 ;
			15'h00003631 : data <= 8'b00000000 ;
			15'h00003632 : data <= 8'b00000000 ;
			15'h00003633 : data <= 8'b00000000 ;
			15'h00003634 : data <= 8'b00000000 ;
			15'h00003635 : data <= 8'b00000000 ;
			15'h00003636 : data <= 8'b00000000 ;
			15'h00003637 : data <= 8'b00000000 ;
			15'h00003638 : data <= 8'b00000000 ;
			15'h00003639 : data <= 8'b00000000 ;
			15'h0000363A : data <= 8'b00000000 ;
			15'h0000363B : data <= 8'b00000000 ;
			15'h0000363C : data <= 8'b00000000 ;
			15'h0000363D : data <= 8'b00000000 ;
			15'h0000363E : data <= 8'b00000000 ;
			15'h0000363F : data <= 8'b00000000 ;
			15'h00003640 : data <= 8'b00000000 ;
			15'h00003641 : data <= 8'b00000000 ;
			15'h00003642 : data <= 8'b00000000 ;
			15'h00003643 : data <= 8'b00000000 ;
			15'h00003644 : data <= 8'b00000000 ;
			15'h00003645 : data <= 8'b00000000 ;
			15'h00003646 : data <= 8'b00000000 ;
			15'h00003647 : data <= 8'b00000000 ;
			15'h00003648 : data <= 8'b00000000 ;
			15'h00003649 : data <= 8'b00000000 ;
			15'h0000364A : data <= 8'b00000000 ;
			15'h0000364B : data <= 8'b00000000 ;
			15'h0000364C : data <= 8'b00000000 ;
			15'h0000364D : data <= 8'b00000000 ;
			15'h0000364E : data <= 8'b00000000 ;
			15'h0000364F : data <= 8'b00000000 ;
			15'h00003650 : data <= 8'b00000000 ;
			15'h00003651 : data <= 8'b00000000 ;
			15'h00003652 : data <= 8'b00000000 ;
			15'h00003653 : data <= 8'b00000000 ;
			15'h00003654 : data <= 8'b00000000 ;
			15'h00003655 : data <= 8'b00000000 ;
			15'h00003656 : data <= 8'b00000000 ;
			15'h00003657 : data <= 8'b00000000 ;
			15'h00003658 : data <= 8'b00000000 ;
			15'h00003659 : data <= 8'b00000000 ;
			15'h0000365A : data <= 8'b00000000 ;
			15'h0000365B : data <= 8'b00000000 ;
			15'h0000365C : data <= 8'b00000000 ;
			15'h0000365D : data <= 8'b00000000 ;
			15'h0000365E : data <= 8'b00000000 ;
			15'h0000365F : data <= 8'b00000000 ;
			15'h00003660 : data <= 8'b00000000 ;
			15'h00003661 : data <= 8'b00000000 ;
			15'h00003662 : data <= 8'b00000000 ;
			15'h00003663 : data <= 8'b00000000 ;
			15'h00003664 : data <= 8'b00000000 ;
			15'h00003665 : data <= 8'b00000000 ;
			15'h00003666 : data <= 8'b00000000 ;
			15'h00003667 : data <= 8'b00000000 ;
			15'h00003668 : data <= 8'b00000000 ;
			15'h00003669 : data <= 8'b00000000 ;
			15'h0000366A : data <= 8'b00000000 ;
			15'h0000366B : data <= 8'b00000000 ;
			15'h0000366C : data <= 8'b00000000 ;
			15'h0000366D : data <= 8'b00000000 ;
			15'h0000366E : data <= 8'b00000000 ;
			15'h0000366F : data <= 8'b00000000 ;
			15'h00003670 : data <= 8'b00000000 ;
			15'h00003671 : data <= 8'b00000000 ;
			15'h00003672 : data <= 8'b00000000 ;
			15'h00003673 : data <= 8'b00000000 ;
			15'h00003674 : data <= 8'b00000000 ;
			15'h00003675 : data <= 8'b00000000 ;
			15'h00003676 : data <= 8'b00000000 ;
			15'h00003677 : data <= 8'b00000000 ;
			15'h00003678 : data <= 8'b00000000 ;
			15'h00003679 : data <= 8'b00000000 ;
			15'h0000367A : data <= 8'b00000000 ;
			15'h0000367B : data <= 8'b00000000 ;
			15'h0000367C : data <= 8'b00000000 ;
			15'h0000367D : data <= 8'b00000000 ;
			15'h0000367E : data <= 8'b00000000 ;
			15'h0000367F : data <= 8'b00000000 ;
			15'h00003680 : data <= 8'b00000000 ;
			15'h00003681 : data <= 8'b00000000 ;
			15'h00003682 : data <= 8'b00000000 ;
			15'h00003683 : data <= 8'b00000000 ;
			15'h00003684 : data <= 8'b00000000 ;
			15'h00003685 : data <= 8'b00000000 ;
			15'h00003686 : data <= 8'b00000000 ;
			15'h00003687 : data <= 8'b00000000 ;
			15'h00003688 : data <= 8'b00000000 ;
			15'h00003689 : data <= 8'b00000000 ;
			15'h0000368A : data <= 8'b00000000 ;
			15'h0000368B : data <= 8'b00000000 ;
			15'h0000368C : data <= 8'b00000000 ;
			15'h0000368D : data <= 8'b00000000 ;
			15'h0000368E : data <= 8'b00000000 ;
			15'h0000368F : data <= 8'b00000000 ;
			15'h00003690 : data <= 8'b00000000 ;
			15'h00003691 : data <= 8'b00000000 ;
			15'h00003692 : data <= 8'b00000000 ;
			15'h00003693 : data <= 8'b00000000 ;
			15'h00003694 : data <= 8'b00000000 ;
			15'h00003695 : data <= 8'b00000000 ;
			15'h00003696 : data <= 8'b00000000 ;
			15'h00003697 : data <= 8'b00000000 ;
			15'h00003698 : data <= 8'b00000000 ;
			15'h00003699 : data <= 8'b00000000 ;
			15'h0000369A : data <= 8'b00000000 ;
			15'h0000369B : data <= 8'b00000000 ;
			15'h0000369C : data <= 8'b00000000 ;
			15'h0000369D : data <= 8'b00000000 ;
			15'h0000369E : data <= 8'b00000000 ;
			15'h0000369F : data <= 8'b00000000 ;
			15'h000036A0 : data <= 8'b00000000 ;
			15'h000036A1 : data <= 8'b00000000 ;
			15'h000036A2 : data <= 8'b00000000 ;
			15'h000036A3 : data <= 8'b00000000 ;
			15'h000036A4 : data <= 8'b00000000 ;
			15'h000036A5 : data <= 8'b00000000 ;
			15'h000036A6 : data <= 8'b00000000 ;
			15'h000036A7 : data <= 8'b00000000 ;
			15'h000036A8 : data <= 8'b00000000 ;
			15'h000036A9 : data <= 8'b00000000 ;
			15'h000036AA : data <= 8'b00000000 ;
			15'h000036AB : data <= 8'b00000000 ;
			15'h000036AC : data <= 8'b00000000 ;
			15'h000036AD : data <= 8'b00000000 ;
			15'h000036AE : data <= 8'b00000000 ;
			15'h000036AF : data <= 8'b00000000 ;
			15'h000036B0 : data <= 8'b00000000 ;
			15'h000036B1 : data <= 8'b00000000 ;
			15'h000036B2 : data <= 8'b00000000 ;
			15'h000036B3 : data <= 8'b00000000 ;
			15'h000036B4 : data <= 8'b00000000 ;
			15'h000036B5 : data <= 8'b00000000 ;
			15'h000036B6 : data <= 8'b00000000 ;
			15'h000036B7 : data <= 8'b00000000 ;
			15'h000036B8 : data <= 8'b00000000 ;
			15'h000036B9 : data <= 8'b00000000 ;
			15'h000036BA : data <= 8'b00000000 ;
			15'h000036BB : data <= 8'b00000000 ;
			15'h000036BC : data <= 8'b00000000 ;
			15'h000036BD : data <= 8'b00000000 ;
			15'h000036BE : data <= 8'b00000000 ;
			15'h000036BF : data <= 8'b00000000 ;
			15'h000036C0 : data <= 8'b00000000 ;
			15'h000036C1 : data <= 8'b00000000 ;
			15'h000036C2 : data <= 8'b00000000 ;
			15'h000036C3 : data <= 8'b00000000 ;
			15'h000036C4 : data <= 8'b00000000 ;
			15'h000036C5 : data <= 8'b00000000 ;
			15'h000036C6 : data <= 8'b00000000 ;
			15'h000036C7 : data <= 8'b00000000 ;
			15'h000036C8 : data <= 8'b00000000 ;
			15'h000036C9 : data <= 8'b00000000 ;
			15'h000036CA : data <= 8'b00000000 ;
			15'h000036CB : data <= 8'b00000000 ;
			15'h000036CC : data <= 8'b00000000 ;
			15'h000036CD : data <= 8'b00000000 ;
			15'h000036CE : data <= 8'b00000000 ;
			15'h000036CF : data <= 8'b00000000 ;
			15'h000036D0 : data <= 8'b00000000 ;
			15'h000036D1 : data <= 8'b00000000 ;
			15'h000036D2 : data <= 8'b00000000 ;
			15'h000036D3 : data <= 8'b00000000 ;
			15'h000036D4 : data <= 8'b00000000 ;
			15'h000036D5 : data <= 8'b00000000 ;
			15'h000036D6 : data <= 8'b00000000 ;
			15'h000036D7 : data <= 8'b00000000 ;
			15'h000036D8 : data <= 8'b00000000 ;
			15'h000036D9 : data <= 8'b00000000 ;
			15'h000036DA : data <= 8'b00000000 ;
			15'h000036DB : data <= 8'b00000000 ;
			15'h000036DC : data <= 8'b00000000 ;
			15'h000036DD : data <= 8'b00000000 ;
			15'h000036DE : data <= 8'b00000000 ;
			15'h000036DF : data <= 8'b00000000 ;
			15'h000036E0 : data <= 8'b00000000 ;
			15'h000036E1 : data <= 8'b00000000 ;
			15'h000036E2 : data <= 8'b00000000 ;
			15'h000036E3 : data <= 8'b00000000 ;
			15'h000036E4 : data <= 8'b00000000 ;
			15'h000036E5 : data <= 8'b00000000 ;
			15'h000036E6 : data <= 8'b00000000 ;
			15'h000036E7 : data <= 8'b00000000 ;
			15'h000036E8 : data <= 8'b00000000 ;
			15'h000036E9 : data <= 8'b00000000 ;
			15'h000036EA : data <= 8'b00000000 ;
			15'h000036EB : data <= 8'b00000000 ;
			15'h000036EC : data <= 8'b00000000 ;
			15'h000036ED : data <= 8'b00000000 ;
			15'h000036EE : data <= 8'b00000000 ;
			15'h000036EF : data <= 8'b00000000 ;
			15'h000036F0 : data <= 8'b00000000 ;
			15'h000036F1 : data <= 8'b00000000 ;
			15'h000036F2 : data <= 8'b00000000 ;
			15'h000036F3 : data <= 8'b00000000 ;
			15'h000036F4 : data <= 8'b00000000 ;
			15'h000036F5 : data <= 8'b00000000 ;
			15'h000036F6 : data <= 8'b00000000 ;
			15'h000036F7 : data <= 8'b00000000 ;
			15'h000036F8 : data <= 8'b00000000 ;
			15'h000036F9 : data <= 8'b00000000 ;
			15'h000036FA : data <= 8'b00000000 ;
			15'h000036FB : data <= 8'b00000000 ;
			15'h000036FC : data <= 8'b00000000 ;
			15'h000036FD : data <= 8'b00000000 ;
			15'h000036FE : data <= 8'b00000000 ;
			15'h000036FF : data <= 8'b00000000 ;
			15'h00003700 : data <= 8'b00000000 ;
			15'h00003701 : data <= 8'b00000000 ;
			15'h00003702 : data <= 8'b00000000 ;
			15'h00003703 : data <= 8'b00000000 ;
			15'h00003704 : data <= 8'b00000000 ;
			15'h00003705 : data <= 8'b00000000 ;
			15'h00003706 : data <= 8'b00000000 ;
			15'h00003707 : data <= 8'b00000000 ;
			15'h00003708 : data <= 8'b00000000 ;
			15'h00003709 : data <= 8'b00000000 ;
			15'h0000370A : data <= 8'b00000000 ;
			15'h0000370B : data <= 8'b00000000 ;
			15'h0000370C : data <= 8'b00000000 ;
			15'h0000370D : data <= 8'b00000000 ;
			15'h0000370E : data <= 8'b00000000 ;
			15'h0000370F : data <= 8'b00000000 ;
			15'h00003710 : data <= 8'b00000000 ;
			15'h00003711 : data <= 8'b00000000 ;
			15'h00003712 : data <= 8'b00000000 ;
			15'h00003713 : data <= 8'b00000000 ;
			15'h00003714 : data <= 8'b00000000 ;
			15'h00003715 : data <= 8'b00000000 ;
			15'h00003716 : data <= 8'b00000000 ;
			15'h00003717 : data <= 8'b00000000 ;
			15'h00003718 : data <= 8'b00000000 ;
			15'h00003719 : data <= 8'b00000000 ;
			15'h0000371A : data <= 8'b00000000 ;
			15'h0000371B : data <= 8'b00000000 ;
			15'h0000371C : data <= 8'b00000000 ;
			15'h0000371D : data <= 8'b00000000 ;
			15'h0000371E : data <= 8'b00000000 ;
			15'h0000371F : data <= 8'b00000000 ;
			15'h00003720 : data <= 8'b00000000 ;
			15'h00003721 : data <= 8'b00000000 ;
			15'h00003722 : data <= 8'b00000000 ;
			15'h00003723 : data <= 8'b00000000 ;
			15'h00003724 : data <= 8'b00000000 ;
			15'h00003725 : data <= 8'b00000000 ;
			15'h00003726 : data <= 8'b00000000 ;
			15'h00003727 : data <= 8'b00000000 ;
			15'h00003728 : data <= 8'b00000000 ;
			15'h00003729 : data <= 8'b00000000 ;
			15'h0000372A : data <= 8'b00000000 ;
			15'h0000372B : data <= 8'b00000000 ;
			15'h0000372C : data <= 8'b00000000 ;
			15'h0000372D : data <= 8'b00000000 ;
			15'h0000372E : data <= 8'b00000000 ;
			15'h0000372F : data <= 8'b00000000 ;
			15'h00003730 : data <= 8'b00000000 ;
			15'h00003731 : data <= 8'b00000000 ;
			15'h00003732 : data <= 8'b00000000 ;
			15'h00003733 : data <= 8'b00000000 ;
			15'h00003734 : data <= 8'b00000000 ;
			15'h00003735 : data <= 8'b00000000 ;
			15'h00003736 : data <= 8'b00000000 ;
			15'h00003737 : data <= 8'b00000000 ;
			15'h00003738 : data <= 8'b00000000 ;
			15'h00003739 : data <= 8'b00000000 ;
			15'h0000373A : data <= 8'b00000000 ;
			15'h0000373B : data <= 8'b00000000 ;
			15'h0000373C : data <= 8'b00000000 ;
			15'h0000373D : data <= 8'b00000000 ;
			15'h0000373E : data <= 8'b00000000 ;
			15'h0000373F : data <= 8'b00000000 ;
			15'h00003740 : data <= 8'b00000000 ;
			15'h00003741 : data <= 8'b00000000 ;
			15'h00003742 : data <= 8'b00000000 ;
			15'h00003743 : data <= 8'b00000000 ;
			15'h00003744 : data <= 8'b00000000 ;
			15'h00003745 : data <= 8'b00000000 ;
			15'h00003746 : data <= 8'b00000000 ;
			15'h00003747 : data <= 8'b00000000 ;
			15'h00003748 : data <= 8'b00000000 ;
			15'h00003749 : data <= 8'b00000000 ;
			15'h0000374A : data <= 8'b00000000 ;
			15'h0000374B : data <= 8'b00000000 ;
			15'h0000374C : data <= 8'b00000000 ;
			15'h0000374D : data <= 8'b00000000 ;
			15'h0000374E : data <= 8'b00000000 ;
			15'h0000374F : data <= 8'b00000000 ;
			15'h00003750 : data <= 8'b00000000 ;
			15'h00003751 : data <= 8'b00000000 ;
			15'h00003752 : data <= 8'b00000000 ;
			15'h00003753 : data <= 8'b00000000 ;
			15'h00003754 : data <= 8'b00000000 ;
			15'h00003755 : data <= 8'b00000000 ;
			15'h00003756 : data <= 8'b00000000 ;
			15'h00003757 : data <= 8'b00000000 ;
			15'h00003758 : data <= 8'b00000000 ;
			15'h00003759 : data <= 8'b00000000 ;
			15'h0000375A : data <= 8'b00000000 ;
			15'h0000375B : data <= 8'b00000000 ;
			15'h0000375C : data <= 8'b00000000 ;
			15'h0000375D : data <= 8'b00000000 ;
			15'h0000375E : data <= 8'b00000000 ;
			15'h0000375F : data <= 8'b00000000 ;
			15'h00003760 : data <= 8'b00000000 ;
			15'h00003761 : data <= 8'b00000000 ;
			15'h00003762 : data <= 8'b00000000 ;
			15'h00003763 : data <= 8'b00000000 ;
			15'h00003764 : data <= 8'b00000000 ;
			15'h00003765 : data <= 8'b00000000 ;
			15'h00003766 : data <= 8'b00000000 ;
			15'h00003767 : data <= 8'b00000000 ;
			15'h00003768 : data <= 8'b00000000 ;
			15'h00003769 : data <= 8'b00000000 ;
			15'h0000376A : data <= 8'b00000000 ;
			15'h0000376B : data <= 8'b00000000 ;
			15'h0000376C : data <= 8'b00000000 ;
			15'h0000376D : data <= 8'b00000000 ;
			15'h0000376E : data <= 8'b00000000 ;
			15'h0000376F : data <= 8'b00000000 ;
			15'h00003770 : data <= 8'b00000000 ;
			15'h00003771 : data <= 8'b00000000 ;
			15'h00003772 : data <= 8'b00000000 ;
			15'h00003773 : data <= 8'b00000000 ;
			15'h00003774 : data <= 8'b00000000 ;
			15'h00003775 : data <= 8'b00000000 ;
			15'h00003776 : data <= 8'b00000000 ;
			15'h00003777 : data <= 8'b00000000 ;
			15'h00003778 : data <= 8'b00000000 ;
			15'h00003779 : data <= 8'b00000000 ;
			15'h0000377A : data <= 8'b00000000 ;
			15'h0000377B : data <= 8'b00000000 ;
			15'h0000377C : data <= 8'b00000000 ;
			15'h0000377D : data <= 8'b00000000 ;
			15'h0000377E : data <= 8'b00000000 ;
			15'h0000377F : data <= 8'b00000000 ;
			15'h00003780 : data <= 8'b00000000 ;
			15'h00003781 : data <= 8'b00000000 ;
			15'h00003782 : data <= 8'b00000000 ;
			15'h00003783 : data <= 8'b00000000 ;
			15'h00003784 : data <= 8'b00000000 ;
			15'h00003785 : data <= 8'b00000000 ;
			15'h00003786 : data <= 8'b00000000 ;
			15'h00003787 : data <= 8'b00000000 ;
			15'h00003788 : data <= 8'b00000000 ;
			15'h00003789 : data <= 8'b00000000 ;
			15'h0000378A : data <= 8'b00000000 ;
			15'h0000378B : data <= 8'b00000000 ;
			15'h0000378C : data <= 8'b00000000 ;
			15'h0000378D : data <= 8'b00000000 ;
			15'h0000378E : data <= 8'b00000000 ;
			15'h0000378F : data <= 8'b00000000 ;
			15'h00003790 : data <= 8'b00000000 ;
			15'h00003791 : data <= 8'b00000000 ;
			15'h00003792 : data <= 8'b00000000 ;
			15'h00003793 : data <= 8'b00000000 ;
			15'h00003794 : data <= 8'b00000000 ;
			15'h00003795 : data <= 8'b00000000 ;
			15'h00003796 : data <= 8'b00000000 ;
			15'h00003797 : data <= 8'b00000000 ;
			15'h00003798 : data <= 8'b00000000 ;
			15'h00003799 : data <= 8'b00000000 ;
			15'h0000379A : data <= 8'b00000000 ;
			15'h0000379B : data <= 8'b00000000 ;
			15'h0000379C : data <= 8'b00000000 ;
			15'h0000379D : data <= 8'b00000000 ;
			15'h0000379E : data <= 8'b00000000 ;
			15'h0000379F : data <= 8'b00000000 ;
			15'h000037A0 : data <= 8'b00000000 ;
			15'h000037A1 : data <= 8'b00000000 ;
			15'h000037A2 : data <= 8'b00000000 ;
			15'h000037A3 : data <= 8'b00000000 ;
			15'h000037A4 : data <= 8'b00000000 ;
			15'h000037A5 : data <= 8'b00000000 ;
			15'h000037A6 : data <= 8'b00000000 ;
			15'h000037A7 : data <= 8'b00000000 ;
			15'h000037A8 : data <= 8'b00000000 ;
			15'h000037A9 : data <= 8'b00000000 ;
			15'h000037AA : data <= 8'b00000000 ;
			15'h000037AB : data <= 8'b00000000 ;
			15'h000037AC : data <= 8'b00000000 ;
			15'h000037AD : data <= 8'b00000000 ;
			15'h000037AE : data <= 8'b00000000 ;
			15'h000037AF : data <= 8'b00000000 ;
			15'h000037B0 : data <= 8'b00000000 ;
			15'h000037B1 : data <= 8'b00000000 ;
			15'h000037B2 : data <= 8'b00000000 ;
			15'h000037B3 : data <= 8'b00000000 ;
			15'h000037B4 : data <= 8'b00000000 ;
			15'h000037B5 : data <= 8'b00000000 ;
			15'h000037B6 : data <= 8'b00000000 ;
			15'h000037B7 : data <= 8'b00000000 ;
			15'h000037B8 : data <= 8'b00000000 ;
			15'h000037B9 : data <= 8'b00000000 ;
			15'h000037BA : data <= 8'b00000000 ;
			15'h000037BB : data <= 8'b00000000 ;
			15'h000037BC : data <= 8'b00000000 ;
			15'h000037BD : data <= 8'b00000000 ;
			15'h000037BE : data <= 8'b00000000 ;
			15'h000037BF : data <= 8'b00000000 ;
			15'h000037C0 : data <= 8'b00000000 ;
			15'h000037C1 : data <= 8'b00000000 ;
			15'h000037C2 : data <= 8'b00000000 ;
			15'h000037C3 : data <= 8'b00000000 ;
			15'h000037C4 : data <= 8'b00000000 ;
			15'h000037C5 : data <= 8'b00000000 ;
			15'h000037C6 : data <= 8'b00000000 ;
			15'h000037C7 : data <= 8'b00000000 ;
			15'h000037C8 : data <= 8'b00000000 ;
			15'h000037C9 : data <= 8'b00000000 ;
			15'h000037CA : data <= 8'b00000000 ;
			15'h000037CB : data <= 8'b00000000 ;
			15'h000037CC : data <= 8'b00000000 ;
			15'h000037CD : data <= 8'b00000000 ;
			15'h000037CE : data <= 8'b00000000 ;
			15'h000037CF : data <= 8'b00000000 ;
			15'h000037D0 : data <= 8'b00000000 ;
			15'h000037D1 : data <= 8'b00000000 ;
			15'h000037D2 : data <= 8'b00000000 ;
			15'h000037D3 : data <= 8'b00000000 ;
			15'h000037D4 : data <= 8'b00000000 ;
			15'h000037D5 : data <= 8'b00000000 ;
			15'h000037D6 : data <= 8'b00000000 ;
			15'h000037D7 : data <= 8'b00000000 ;
			15'h000037D8 : data <= 8'b00000000 ;
			15'h000037D9 : data <= 8'b00000000 ;
			15'h000037DA : data <= 8'b00000000 ;
			15'h000037DB : data <= 8'b00000000 ;
			15'h000037DC : data <= 8'b00000000 ;
			15'h000037DD : data <= 8'b00000000 ;
			15'h000037DE : data <= 8'b00000000 ;
			15'h000037DF : data <= 8'b00000000 ;
			15'h000037E0 : data <= 8'b00000000 ;
			15'h000037E1 : data <= 8'b00000000 ;
			15'h000037E2 : data <= 8'b00000000 ;
			15'h000037E3 : data <= 8'b00000000 ;
			15'h000037E4 : data <= 8'b00000000 ;
			15'h000037E5 : data <= 8'b00000000 ;
			15'h000037E6 : data <= 8'b00000000 ;
			15'h000037E7 : data <= 8'b00000000 ;
			15'h000037E8 : data <= 8'b00000000 ;
			15'h000037E9 : data <= 8'b00000000 ;
			15'h000037EA : data <= 8'b00000000 ;
			15'h000037EB : data <= 8'b00000000 ;
			15'h000037EC : data <= 8'b00000000 ;
			15'h000037ED : data <= 8'b00000000 ;
			15'h000037EE : data <= 8'b00000000 ;
			15'h000037EF : data <= 8'b00000000 ;
			15'h000037F0 : data <= 8'b00000000 ;
			15'h000037F1 : data <= 8'b00000000 ;
			15'h000037F2 : data <= 8'b00000000 ;
			15'h000037F3 : data <= 8'b00000000 ;
			15'h000037F4 : data <= 8'b00000000 ;
			15'h000037F5 : data <= 8'b00000000 ;
			15'h000037F6 : data <= 8'b00000000 ;
			15'h000037F7 : data <= 8'b00000000 ;
			15'h000037F8 : data <= 8'b00000000 ;
			15'h000037F9 : data <= 8'b00000000 ;
			15'h000037FA : data <= 8'b00000000 ;
			15'h000037FB : data <= 8'b00000000 ;
			15'h000037FC : data <= 8'b00000000 ;
			15'h000037FD : data <= 8'b00000000 ;
			15'h000037FE : data <= 8'b00000000 ;
			15'h000037FF : data <= 8'b00000000 ;
			15'h00003800 : data <= 8'b00000000 ;
			15'h00003801 : data <= 8'b00000000 ;
			15'h00003802 : data <= 8'b00000000 ;
			15'h00003803 : data <= 8'b00000000 ;
			15'h00003804 : data <= 8'b00000000 ;
			15'h00003805 : data <= 8'b00000000 ;
			15'h00003806 : data <= 8'b00000000 ;
			15'h00003807 : data <= 8'b00000000 ;
			15'h00003808 : data <= 8'b00000000 ;
			15'h00003809 : data <= 8'b00000000 ;
			15'h0000380A : data <= 8'b00000000 ;
			15'h0000380B : data <= 8'b00000000 ;
			15'h0000380C : data <= 8'b00000000 ;
			15'h0000380D : data <= 8'b00000000 ;
			15'h0000380E : data <= 8'b00000000 ;
			15'h0000380F : data <= 8'b00000000 ;
			15'h00003810 : data <= 8'b00000000 ;
			15'h00003811 : data <= 8'b00000000 ;
			15'h00003812 : data <= 8'b00000000 ;
			15'h00003813 : data <= 8'b00000000 ;
			15'h00003814 : data <= 8'b00000000 ;
			15'h00003815 : data <= 8'b00000000 ;
			15'h00003816 : data <= 8'b00000000 ;
			15'h00003817 : data <= 8'b00000000 ;
			15'h00003818 : data <= 8'b00000000 ;
			15'h00003819 : data <= 8'b00000000 ;
			15'h0000381A : data <= 8'b00000000 ;
			15'h0000381B : data <= 8'b00000000 ;
			15'h0000381C : data <= 8'b00000000 ;
			15'h0000381D : data <= 8'b00000000 ;
			15'h0000381E : data <= 8'b00000000 ;
			15'h0000381F : data <= 8'b00000000 ;
			15'h00003820 : data <= 8'b00000000 ;
			15'h00003821 : data <= 8'b00000000 ;
			15'h00003822 : data <= 8'b00000000 ;
			15'h00003823 : data <= 8'b00000000 ;
			15'h00003824 : data <= 8'b00000000 ;
			15'h00003825 : data <= 8'b00000000 ;
			15'h00003826 : data <= 8'b00000000 ;
			15'h00003827 : data <= 8'b00000000 ;
			15'h00003828 : data <= 8'b00000000 ;
			15'h00003829 : data <= 8'b00000000 ;
			15'h0000382A : data <= 8'b00000000 ;
			15'h0000382B : data <= 8'b00000000 ;
			15'h0000382C : data <= 8'b00000000 ;
			15'h0000382D : data <= 8'b00000000 ;
			15'h0000382E : data <= 8'b00000000 ;
			15'h0000382F : data <= 8'b00000000 ;
			15'h00003830 : data <= 8'b00000000 ;
			15'h00003831 : data <= 8'b00000000 ;
			15'h00003832 : data <= 8'b00000000 ;
			15'h00003833 : data <= 8'b00000000 ;
			15'h00003834 : data <= 8'b00000000 ;
			15'h00003835 : data <= 8'b00000000 ;
			15'h00003836 : data <= 8'b00000000 ;
			15'h00003837 : data <= 8'b00000000 ;
			15'h00003838 : data <= 8'b00000000 ;
			15'h00003839 : data <= 8'b00000000 ;
			15'h0000383A : data <= 8'b00000000 ;
			15'h0000383B : data <= 8'b00000000 ;
			15'h0000383C : data <= 8'b00000000 ;
			15'h0000383D : data <= 8'b00000000 ;
			15'h0000383E : data <= 8'b00000000 ;
			15'h0000383F : data <= 8'b00000000 ;
			15'h00003840 : data <= 8'b00000000 ;
			15'h00003841 : data <= 8'b00000000 ;
			15'h00003842 : data <= 8'b00000000 ;
			15'h00003843 : data <= 8'b00000000 ;
			15'h00003844 : data <= 8'b00000000 ;
			15'h00003845 : data <= 8'b00000000 ;
			15'h00003846 : data <= 8'b00000000 ;
			15'h00003847 : data <= 8'b00000000 ;
			15'h00003848 : data <= 8'b00000000 ;
			15'h00003849 : data <= 8'b00000000 ;
			15'h0000384A : data <= 8'b00000000 ;
			15'h0000384B : data <= 8'b00000000 ;
			15'h0000384C : data <= 8'b00000000 ;
			15'h0000384D : data <= 8'b00000000 ;
			15'h0000384E : data <= 8'b00000000 ;
			15'h0000384F : data <= 8'b00000000 ;
			15'h00003850 : data <= 8'b00000000 ;
			15'h00003851 : data <= 8'b00000000 ;
			15'h00003852 : data <= 8'b00000000 ;
			15'h00003853 : data <= 8'b00000000 ;
			15'h00003854 : data <= 8'b00000000 ;
			15'h00003855 : data <= 8'b00000000 ;
			15'h00003856 : data <= 8'b00000000 ;
			15'h00003857 : data <= 8'b00000000 ;
			15'h00003858 : data <= 8'b00000000 ;
			15'h00003859 : data <= 8'b00000000 ;
			15'h0000385A : data <= 8'b00000000 ;
			15'h0000385B : data <= 8'b00000000 ;
			15'h0000385C : data <= 8'b00000000 ;
			15'h0000385D : data <= 8'b00000000 ;
			15'h0000385E : data <= 8'b00000000 ;
			15'h0000385F : data <= 8'b00000000 ;
			15'h00003860 : data <= 8'b00000000 ;
			15'h00003861 : data <= 8'b00000000 ;
			15'h00003862 : data <= 8'b00000000 ;
			15'h00003863 : data <= 8'b00000000 ;
			15'h00003864 : data <= 8'b00000000 ;
			15'h00003865 : data <= 8'b00000000 ;
			15'h00003866 : data <= 8'b00000000 ;
			15'h00003867 : data <= 8'b00000000 ;
			15'h00003868 : data <= 8'b00000000 ;
			15'h00003869 : data <= 8'b00000000 ;
			15'h0000386A : data <= 8'b00000000 ;
			15'h0000386B : data <= 8'b00000000 ;
			15'h0000386C : data <= 8'b00000000 ;
			15'h0000386D : data <= 8'b00000000 ;
			15'h0000386E : data <= 8'b00000000 ;
			15'h0000386F : data <= 8'b00000000 ;
			15'h00003870 : data <= 8'b00000000 ;
			15'h00003871 : data <= 8'b00000000 ;
			15'h00003872 : data <= 8'b00000000 ;
			15'h00003873 : data <= 8'b00000000 ;
			15'h00003874 : data <= 8'b00000000 ;
			15'h00003875 : data <= 8'b00000000 ;
			15'h00003876 : data <= 8'b00000000 ;
			15'h00003877 : data <= 8'b00000000 ;
			15'h00003878 : data <= 8'b00000000 ;
			15'h00003879 : data <= 8'b00000000 ;
			15'h0000387A : data <= 8'b00000000 ;
			15'h0000387B : data <= 8'b00000000 ;
			15'h0000387C : data <= 8'b00000000 ;
			15'h0000387D : data <= 8'b00000000 ;
			15'h0000387E : data <= 8'b00000000 ;
			15'h0000387F : data <= 8'b00000000 ;
			15'h00003880 : data <= 8'b00000000 ;
			15'h00003881 : data <= 8'b00000000 ;
			15'h00003882 : data <= 8'b00000000 ;
			15'h00003883 : data <= 8'b00000000 ;
			15'h00003884 : data <= 8'b00000000 ;
			15'h00003885 : data <= 8'b00000000 ;
			15'h00003886 : data <= 8'b00000000 ;
			15'h00003887 : data <= 8'b00000000 ;
			15'h00003888 : data <= 8'b00000000 ;
			15'h00003889 : data <= 8'b00000000 ;
			15'h0000388A : data <= 8'b00000000 ;
			15'h0000388B : data <= 8'b00000000 ;
			15'h0000388C : data <= 8'b00000000 ;
			15'h0000388D : data <= 8'b00000000 ;
			15'h0000388E : data <= 8'b00000000 ;
			15'h0000388F : data <= 8'b00000000 ;
			15'h00003890 : data <= 8'b00000000 ;
			15'h00003891 : data <= 8'b00000000 ;
			15'h00003892 : data <= 8'b00000000 ;
			15'h00003893 : data <= 8'b00000000 ;
			15'h00003894 : data <= 8'b00000000 ;
			15'h00003895 : data <= 8'b00000000 ;
			15'h00003896 : data <= 8'b00000000 ;
			15'h00003897 : data <= 8'b00000000 ;
			15'h00003898 : data <= 8'b00000000 ;
			15'h00003899 : data <= 8'b00000000 ;
			15'h0000389A : data <= 8'b00000000 ;
			15'h0000389B : data <= 8'b00000000 ;
			15'h0000389C : data <= 8'b00000000 ;
			15'h0000389D : data <= 8'b00000000 ;
			15'h0000389E : data <= 8'b00000000 ;
			15'h0000389F : data <= 8'b00000000 ;
			15'h000038A0 : data <= 8'b00000000 ;
			15'h000038A1 : data <= 8'b00000000 ;
			15'h000038A2 : data <= 8'b00000000 ;
			15'h000038A3 : data <= 8'b00000000 ;
			15'h000038A4 : data <= 8'b00000000 ;
			15'h000038A5 : data <= 8'b00000000 ;
			15'h000038A6 : data <= 8'b00000000 ;
			15'h000038A7 : data <= 8'b00000000 ;
			15'h000038A8 : data <= 8'b00000000 ;
			15'h000038A9 : data <= 8'b00000000 ;
			15'h000038AA : data <= 8'b00000000 ;
			15'h000038AB : data <= 8'b00000000 ;
			15'h000038AC : data <= 8'b00000000 ;
			15'h000038AD : data <= 8'b00000000 ;
			15'h000038AE : data <= 8'b00000000 ;
			15'h000038AF : data <= 8'b00000000 ;
			15'h000038B0 : data <= 8'b00000000 ;
			15'h000038B1 : data <= 8'b00000000 ;
			15'h000038B2 : data <= 8'b00000000 ;
			15'h000038B3 : data <= 8'b00000000 ;
			15'h000038B4 : data <= 8'b00000000 ;
			15'h000038B5 : data <= 8'b00000000 ;
			15'h000038B6 : data <= 8'b00000000 ;
			15'h000038B7 : data <= 8'b00000000 ;
			15'h000038B8 : data <= 8'b00000000 ;
			15'h000038B9 : data <= 8'b00000000 ;
			15'h000038BA : data <= 8'b00000000 ;
			15'h000038BB : data <= 8'b00000000 ;
			15'h000038BC : data <= 8'b00000000 ;
			15'h000038BD : data <= 8'b00000000 ;
			15'h000038BE : data <= 8'b00000000 ;
			15'h000038BF : data <= 8'b00000000 ;
			15'h000038C0 : data <= 8'b00000000 ;
			15'h000038C1 : data <= 8'b00000000 ;
			15'h000038C2 : data <= 8'b00000000 ;
			15'h000038C3 : data <= 8'b00000000 ;
			15'h000038C4 : data <= 8'b00000000 ;
			15'h000038C5 : data <= 8'b00000000 ;
			15'h000038C6 : data <= 8'b00000000 ;
			15'h000038C7 : data <= 8'b00000000 ;
			15'h000038C8 : data <= 8'b00000000 ;
			15'h000038C9 : data <= 8'b00000000 ;
			15'h000038CA : data <= 8'b00000000 ;
			15'h000038CB : data <= 8'b00000000 ;
			15'h000038CC : data <= 8'b00000000 ;
			15'h000038CD : data <= 8'b00000000 ;
			15'h000038CE : data <= 8'b00000000 ;
			15'h000038CF : data <= 8'b00000000 ;
			15'h000038D0 : data <= 8'b00000000 ;
			15'h000038D1 : data <= 8'b00000000 ;
			15'h000038D2 : data <= 8'b00000000 ;
			15'h000038D3 : data <= 8'b00000000 ;
			15'h000038D4 : data <= 8'b00000000 ;
			15'h000038D5 : data <= 8'b00000000 ;
			15'h000038D6 : data <= 8'b00000000 ;
			15'h000038D7 : data <= 8'b00000000 ;
			15'h000038D8 : data <= 8'b00000000 ;
			15'h000038D9 : data <= 8'b00000000 ;
			15'h000038DA : data <= 8'b00000000 ;
			15'h000038DB : data <= 8'b00000000 ;
			15'h000038DC : data <= 8'b00000000 ;
			15'h000038DD : data <= 8'b00000000 ;
			15'h000038DE : data <= 8'b00000000 ;
			15'h000038DF : data <= 8'b00000000 ;
			15'h000038E0 : data <= 8'b00000000 ;
			15'h000038E1 : data <= 8'b00000000 ;
			15'h000038E2 : data <= 8'b00000000 ;
			15'h000038E3 : data <= 8'b00000000 ;
			15'h000038E4 : data <= 8'b00000000 ;
			15'h000038E5 : data <= 8'b00000000 ;
			15'h000038E6 : data <= 8'b00000000 ;
			15'h000038E7 : data <= 8'b00000000 ;
			15'h000038E8 : data <= 8'b00000000 ;
			15'h000038E9 : data <= 8'b00000000 ;
			15'h000038EA : data <= 8'b00000000 ;
			15'h000038EB : data <= 8'b00000000 ;
			15'h000038EC : data <= 8'b00000000 ;
			15'h000038ED : data <= 8'b00000000 ;
			15'h000038EE : data <= 8'b00000000 ;
			15'h000038EF : data <= 8'b00000000 ;
			15'h000038F0 : data <= 8'b00000000 ;
			15'h000038F1 : data <= 8'b00000000 ;
			15'h000038F2 : data <= 8'b00000000 ;
			15'h000038F3 : data <= 8'b00000000 ;
			15'h000038F4 : data <= 8'b00000000 ;
			15'h000038F5 : data <= 8'b00000000 ;
			15'h000038F6 : data <= 8'b00000000 ;
			15'h000038F7 : data <= 8'b00000000 ;
			15'h000038F8 : data <= 8'b00000000 ;
			15'h000038F9 : data <= 8'b00000000 ;
			15'h000038FA : data <= 8'b00000000 ;
			15'h000038FB : data <= 8'b00000000 ;
			15'h000038FC : data <= 8'b00000000 ;
			15'h000038FD : data <= 8'b00000000 ;
			15'h000038FE : data <= 8'b00000000 ;
			15'h000038FF : data <= 8'b00000000 ;
			15'h00003900 : data <= 8'b00000000 ;
			15'h00003901 : data <= 8'b00000000 ;
			15'h00003902 : data <= 8'b00000000 ;
			15'h00003903 : data <= 8'b00000000 ;
			15'h00003904 : data <= 8'b00000000 ;
			15'h00003905 : data <= 8'b00000000 ;
			15'h00003906 : data <= 8'b00000000 ;
			15'h00003907 : data <= 8'b00000000 ;
			15'h00003908 : data <= 8'b00000000 ;
			15'h00003909 : data <= 8'b00000000 ;
			15'h0000390A : data <= 8'b00000000 ;
			15'h0000390B : data <= 8'b00000000 ;
			15'h0000390C : data <= 8'b00000000 ;
			15'h0000390D : data <= 8'b00000000 ;
			15'h0000390E : data <= 8'b00000000 ;
			15'h0000390F : data <= 8'b00000000 ;
			15'h00003910 : data <= 8'b00000000 ;
			15'h00003911 : data <= 8'b00000000 ;
			15'h00003912 : data <= 8'b00000000 ;
			15'h00003913 : data <= 8'b00000000 ;
			15'h00003914 : data <= 8'b00000000 ;
			15'h00003915 : data <= 8'b00000000 ;
			15'h00003916 : data <= 8'b00000000 ;
			15'h00003917 : data <= 8'b00000000 ;
			15'h00003918 : data <= 8'b00000000 ;
			15'h00003919 : data <= 8'b00000000 ;
			15'h0000391A : data <= 8'b00000000 ;
			15'h0000391B : data <= 8'b00000000 ;
			15'h0000391C : data <= 8'b00000000 ;
			15'h0000391D : data <= 8'b00000000 ;
			15'h0000391E : data <= 8'b00000000 ;
			15'h0000391F : data <= 8'b00000000 ;
			15'h00003920 : data <= 8'b00000000 ;
			15'h00003921 : data <= 8'b00000000 ;
			15'h00003922 : data <= 8'b00000000 ;
			15'h00003923 : data <= 8'b00000000 ;
			15'h00003924 : data <= 8'b00000000 ;
			15'h00003925 : data <= 8'b00000000 ;
			15'h00003926 : data <= 8'b00000000 ;
			15'h00003927 : data <= 8'b00000000 ;
			15'h00003928 : data <= 8'b00000000 ;
			15'h00003929 : data <= 8'b00000000 ;
			15'h0000392A : data <= 8'b00000000 ;
			15'h0000392B : data <= 8'b00000000 ;
			15'h0000392C : data <= 8'b00000000 ;
			15'h0000392D : data <= 8'b00000000 ;
			15'h0000392E : data <= 8'b00000000 ;
			15'h0000392F : data <= 8'b00000000 ;
			15'h00003930 : data <= 8'b00000000 ;
			15'h00003931 : data <= 8'b00000000 ;
			15'h00003932 : data <= 8'b00000000 ;
			15'h00003933 : data <= 8'b00000000 ;
			15'h00003934 : data <= 8'b00000000 ;
			15'h00003935 : data <= 8'b00000000 ;
			15'h00003936 : data <= 8'b00000000 ;
			15'h00003937 : data <= 8'b00000000 ;
			15'h00003938 : data <= 8'b00000000 ;
			15'h00003939 : data <= 8'b00000000 ;
			15'h0000393A : data <= 8'b00000000 ;
			15'h0000393B : data <= 8'b00000000 ;
			15'h0000393C : data <= 8'b00000000 ;
			15'h0000393D : data <= 8'b00000000 ;
			15'h0000393E : data <= 8'b00000000 ;
			15'h0000393F : data <= 8'b00000000 ;
			15'h00003940 : data <= 8'b00000000 ;
			15'h00003941 : data <= 8'b00000000 ;
			15'h00003942 : data <= 8'b00000000 ;
			15'h00003943 : data <= 8'b00000000 ;
			15'h00003944 : data <= 8'b00000000 ;
			15'h00003945 : data <= 8'b00000000 ;
			15'h00003946 : data <= 8'b00000000 ;
			15'h00003947 : data <= 8'b00000000 ;
			15'h00003948 : data <= 8'b00000000 ;
			15'h00003949 : data <= 8'b00000000 ;
			15'h0000394A : data <= 8'b00000000 ;
			15'h0000394B : data <= 8'b00000000 ;
			15'h0000394C : data <= 8'b00000000 ;
			15'h0000394D : data <= 8'b00000000 ;
			15'h0000394E : data <= 8'b00000000 ;
			15'h0000394F : data <= 8'b00000000 ;
			15'h00003950 : data <= 8'b00000000 ;
			15'h00003951 : data <= 8'b00000000 ;
			15'h00003952 : data <= 8'b00000000 ;
			15'h00003953 : data <= 8'b00000000 ;
			15'h00003954 : data <= 8'b00000000 ;
			15'h00003955 : data <= 8'b00000000 ;
			15'h00003956 : data <= 8'b00000000 ;
			15'h00003957 : data <= 8'b00000000 ;
			15'h00003958 : data <= 8'b00000000 ;
			15'h00003959 : data <= 8'b00000000 ;
			15'h0000395A : data <= 8'b00000000 ;
			15'h0000395B : data <= 8'b00000000 ;
			15'h0000395C : data <= 8'b00000000 ;
			15'h0000395D : data <= 8'b00000000 ;
			15'h0000395E : data <= 8'b00000000 ;
			15'h0000395F : data <= 8'b00000000 ;
			15'h00003960 : data <= 8'b00000000 ;
			15'h00003961 : data <= 8'b00000000 ;
			15'h00003962 : data <= 8'b00000000 ;
			15'h00003963 : data <= 8'b00000000 ;
			15'h00003964 : data <= 8'b00000000 ;
			15'h00003965 : data <= 8'b00000000 ;
			15'h00003966 : data <= 8'b00000000 ;
			15'h00003967 : data <= 8'b00000000 ;
			15'h00003968 : data <= 8'b00000000 ;
			15'h00003969 : data <= 8'b00000000 ;
			15'h0000396A : data <= 8'b00000000 ;
			15'h0000396B : data <= 8'b00000000 ;
			15'h0000396C : data <= 8'b00000000 ;
			15'h0000396D : data <= 8'b00000000 ;
			15'h0000396E : data <= 8'b00000000 ;
			15'h0000396F : data <= 8'b00000000 ;
			15'h00003970 : data <= 8'b00000000 ;
			15'h00003971 : data <= 8'b00000000 ;
			15'h00003972 : data <= 8'b00000000 ;
			15'h00003973 : data <= 8'b00000000 ;
			15'h00003974 : data <= 8'b00000000 ;
			15'h00003975 : data <= 8'b00000000 ;
			15'h00003976 : data <= 8'b00000000 ;
			15'h00003977 : data <= 8'b00000000 ;
			15'h00003978 : data <= 8'b00000000 ;
			15'h00003979 : data <= 8'b00000000 ;
			15'h0000397A : data <= 8'b00000000 ;
			15'h0000397B : data <= 8'b00000000 ;
			15'h0000397C : data <= 8'b00000000 ;
			15'h0000397D : data <= 8'b00000000 ;
			15'h0000397E : data <= 8'b00000000 ;
			15'h0000397F : data <= 8'b00000000 ;
			15'h00003980 : data <= 8'b00000000 ;
			15'h00003981 : data <= 8'b00000000 ;
			15'h00003982 : data <= 8'b00000000 ;
			15'h00003983 : data <= 8'b00000000 ;
			15'h00003984 : data <= 8'b00000000 ;
			15'h00003985 : data <= 8'b00000000 ;
			15'h00003986 : data <= 8'b00000000 ;
			15'h00003987 : data <= 8'b00000000 ;
			15'h00003988 : data <= 8'b00000000 ;
			15'h00003989 : data <= 8'b00000000 ;
			15'h0000398A : data <= 8'b00000000 ;
			15'h0000398B : data <= 8'b00000000 ;
			15'h0000398C : data <= 8'b00000000 ;
			15'h0000398D : data <= 8'b00000000 ;
			15'h0000398E : data <= 8'b00000000 ;
			15'h0000398F : data <= 8'b00000000 ;
			15'h00003990 : data <= 8'b00000000 ;
			15'h00003991 : data <= 8'b00000000 ;
			15'h00003992 : data <= 8'b00000000 ;
			15'h00003993 : data <= 8'b00000000 ;
			15'h00003994 : data <= 8'b00000000 ;
			15'h00003995 : data <= 8'b00000000 ;
			15'h00003996 : data <= 8'b00000000 ;
			15'h00003997 : data <= 8'b00000000 ;
			15'h00003998 : data <= 8'b00000000 ;
			15'h00003999 : data <= 8'b00000000 ;
			15'h0000399A : data <= 8'b00000000 ;
			15'h0000399B : data <= 8'b00000000 ;
			15'h0000399C : data <= 8'b00000000 ;
			15'h0000399D : data <= 8'b00000000 ;
			15'h0000399E : data <= 8'b00000000 ;
			15'h0000399F : data <= 8'b00000000 ;
			15'h000039A0 : data <= 8'b00000000 ;
			15'h000039A1 : data <= 8'b00000000 ;
			15'h000039A2 : data <= 8'b00000000 ;
			15'h000039A3 : data <= 8'b00000000 ;
			15'h000039A4 : data <= 8'b00000000 ;
			15'h000039A5 : data <= 8'b00000000 ;
			15'h000039A6 : data <= 8'b00000000 ;
			15'h000039A7 : data <= 8'b00000000 ;
			15'h000039A8 : data <= 8'b00000000 ;
			15'h000039A9 : data <= 8'b00000000 ;
			15'h000039AA : data <= 8'b00000000 ;
			15'h000039AB : data <= 8'b00000000 ;
			15'h000039AC : data <= 8'b00000000 ;
			15'h000039AD : data <= 8'b00000000 ;
			15'h000039AE : data <= 8'b00000000 ;
			15'h000039AF : data <= 8'b00000000 ;
			15'h000039B0 : data <= 8'b00000000 ;
			15'h000039B1 : data <= 8'b00000000 ;
			15'h000039B2 : data <= 8'b00000000 ;
			15'h000039B3 : data <= 8'b00000000 ;
			15'h000039B4 : data <= 8'b00000000 ;
			15'h000039B5 : data <= 8'b00000000 ;
			15'h000039B6 : data <= 8'b00000000 ;
			15'h000039B7 : data <= 8'b00000000 ;
			15'h000039B8 : data <= 8'b00000000 ;
			15'h000039B9 : data <= 8'b00000000 ;
			15'h000039BA : data <= 8'b00000000 ;
			15'h000039BB : data <= 8'b00000000 ;
			15'h000039BC : data <= 8'b00000000 ;
			15'h000039BD : data <= 8'b00000000 ;
			15'h000039BE : data <= 8'b00000000 ;
			15'h000039BF : data <= 8'b00000000 ;
			15'h000039C0 : data <= 8'b00000000 ;
			15'h000039C1 : data <= 8'b00000000 ;
			15'h000039C2 : data <= 8'b00000000 ;
			15'h000039C3 : data <= 8'b00000000 ;
			15'h000039C4 : data <= 8'b00000000 ;
			15'h000039C5 : data <= 8'b00000000 ;
			15'h000039C6 : data <= 8'b00000000 ;
			15'h000039C7 : data <= 8'b00000000 ;
			15'h000039C8 : data <= 8'b00000000 ;
			15'h000039C9 : data <= 8'b00000000 ;
			15'h000039CA : data <= 8'b00000000 ;
			15'h000039CB : data <= 8'b00000000 ;
			15'h000039CC : data <= 8'b00000000 ;
			15'h000039CD : data <= 8'b00000000 ;
			15'h000039CE : data <= 8'b00000000 ;
			15'h000039CF : data <= 8'b00000000 ;
			15'h000039D0 : data <= 8'b00000000 ;
			15'h000039D1 : data <= 8'b00000000 ;
			15'h000039D2 : data <= 8'b00000000 ;
			15'h000039D3 : data <= 8'b00000000 ;
			15'h000039D4 : data <= 8'b00000000 ;
			15'h000039D5 : data <= 8'b00000000 ;
			15'h000039D6 : data <= 8'b00000000 ;
			15'h000039D7 : data <= 8'b00000000 ;
			15'h000039D8 : data <= 8'b00000000 ;
			15'h000039D9 : data <= 8'b00000000 ;
			15'h000039DA : data <= 8'b00000000 ;
			15'h000039DB : data <= 8'b00000000 ;
			15'h000039DC : data <= 8'b00000000 ;
			15'h000039DD : data <= 8'b00000000 ;
			15'h000039DE : data <= 8'b00000000 ;
			15'h000039DF : data <= 8'b00000000 ;
			15'h000039E0 : data <= 8'b00000000 ;
			15'h000039E1 : data <= 8'b00000000 ;
			15'h000039E2 : data <= 8'b00000000 ;
			15'h000039E3 : data <= 8'b00000000 ;
			15'h000039E4 : data <= 8'b00000000 ;
			15'h000039E5 : data <= 8'b00000000 ;
			15'h000039E6 : data <= 8'b00000000 ;
			15'h000039E7 : data <= 8'b00000000 ;
			15'h000039E8 : data <= 8'b00000000 ;
			15'h000039E9 : data <= 8'b00000000 ;
			15'h000039EA : data <= 8'b00000000 ;
			15'h000039EB : data <= 8'b00000000 ;
			15'h000039EC : data <= 8'b00000000 ;
			15'h000039ED : data <= 8'b00000000 ;
			15'h000039EE : data <= 8'b00000000 ;
			15'h000039EF : data <= 8'b00000000 ;
			15'h000039F0 : data <= 8'b00000000 ;
			15'h000039F1 : data <= 8'b00000000 ;
			15'h000039F2 : data <= 8'b00000000 ;
			15'h000039F3 : data <= 8'b00000000 ;
			15'h000039F4 : data <= 8'b00000000 ;
			15'h000039F5 : data <= 8'b00000000 ;
			15'h000039F6 : data <= 8'b00000000 ;
			15'h000039F7 : data <= 8'b00000000 ;
			15'h000039F8 : data <= 8'b00000000 ;
			15'h000039F9 : data <= 8'b00000000 ;
			15'h000039FA : data <= 8'b00000000 ;
			15'h000039FB : data <= 8'b00000000 ;
			15'h000039FC : data <= 8'b00000000 ;
			15'h000039FD : data <= 8'b00000000 ;
			15'h000039FE : data <= 8'b00000000 ;
			15'h000039FF : data <= 8'b00000000 ;
			15'h00003A00 : data <= 8'b00000000 ;
			15'h00003A01 : data <= 8'b00000000 ;
			15'h00003A02 : data <= 8'b00000000 ;
			15'h00003A03 : data <= 8'b00000000 ;
			15'h00003A04 : data <= 8'b00000000 ;
			15'h00003A05 : data <= 8'b00000000 ;
			15'h00003A06 : data <= 8'b00000000 ;
			15'h00003A07 : data <= 8'b00000000 ;
			15'h00003A08 : data <= 8'b00000000 ;
			15'h00003A09 : data <= 8'b00000000 ;
			15'h00003A0A : data <= 8'b00000000 ;
			15'h00003A0B : data <= 8'b00000000 ;
			15'h00003A0C : data <= 8'b00000000 ;
			15'h00003A0D : data <= 8'b00000000 ;
			15'h00003A0E : data <= 8'b00000000 ;
			15'h00003A0F : data <= 8'b00000000 ;
			15'h00003A10 : data <= 8'b00000000 ;
			15'h00003A11 : data <= 8'b00000000 ;
			15'h00003A12 : data <= 8'b00000000 ;
			15'h00003A13 : data <= 8'b00000000 ;
			15'h00003A14 : data <= 8'b00000000 ;
			15'h00003A15 : data <= 8'b00000000 ;
			15'h00003A16 : data <= 8'b00000000 ;
			15'h00003A17 : data <= 8'b00000000 ;
			15'h00003A18 : data <= 8'b00000000 ;
			15'h00003A19 : data <= 8'b00000000 ;
			15'h00003A1A : data <= 8'b00000000 ;
			15'h00003A1B : data <= 8'b00000000 ;
			15'h00003A1C : data <= 8'b00000000 ;
			15'h00003A1D : data <= 8'b00000000 ;
			15'h00003A1E : data <= 8'b00000000 ;
			15'h00003A1F : data <= 8'b00000000 ;
			15'h00003A20 : data <= 8'b00000000 ;
			15'h00003A21 : data <= 8'b00000000 ;
			15'h00003A22 : data <= 8'b00000000 ;
			15'h00003A23 : data <= 8'b00000000 ;
			15'h00003A24 : data <= 8'b00000000 ;
			15'h00003A25 : data <= 8'b00000000 ;
			15'h00003A26 : data <= 8'b00000000 ;
			15'h00003A27 : data <= 8'b00000000 ;
			15'h00003A28 : data <= 8'b00000000 ;
			15'h00003A29 : data <= 8'b00000000 ;
			15'h00003A2A : data <= 8'b00000000 ;
			15'h00003A2B : data <= 8'b00000000 ;
			15'h00003A2C : data <= 8'b00000000 ;
			15'h00003A2D : data <= 8'b00000000 ;
			15'h00003A2E : data <= 8'b00000000 ;
			15'h00003A2F : data <= 8'b00000000 ;
			15'h00003A30 : data <= 8'b00000000 ;
			15'h00003A31 : data <= 8'b00000000 ;
			15'h00003A32 : data <= 8'b00000000 ;
			15'h00003A33 : data <= 8'b00000000 ;
			15'h00003A34 : data <= 8'b00000000 ;
			15'h00003A35 : data <= 8'b00000000 ;
			15'h00003A36 : data <= 8'b00000000 ;
			15'h00003A37 : data <= 8'b00000000 ;
			15'h00003A38 : data <= 8'b00000000 ;
			15'h00003A39 : data <= 8'b00000000 ;
			15'h00003A3A : data <= 8'b00000000 ;
			15'h00003A3B : data <= 8'b00000000 ;
			15'h00003A3C : data <= 8'b00000000 ;
			15'h00003A3D : data <= 8'b00000000 ;
			15'h00003A3E : data <= 8'b00000000 ;
			15'h00003A3F : data <= 8'b00000000 ;
			15'h00003A40 : data <= 8'b00000000 ;
			15'h00003A41 : data <= 8'b00000000 ;
			15'h00003A42 : data <= 8'b00000000 ;
			15'h00003A43 : data <= 8'b00000000 ;
			15'h00003A44 : data <= 8'b00000000 ;
			15'h00003A45 : data <= 8'b00000000 ;
			15'h00003A46 : data <= 8'b00000000 ;
			15'h00003A47 : data <= 8'b00000000 ;
			15'h00003A48 : data <= 8'b00000000 ;
			15'h00003A49 : data <= 8'b00000000 ;
			15'h00003A4A : data <= 8'b00000000 ;
			15'h00003A4B : data <= 8'b00000000 ;
			15'h00003A4C : data <= 8'b00000000 ;
			15'h00003A4D : data <= 8'b00000000 ;
			15'h00003A4E : data <= 8'b00000000 ;
			15'h00003A4F : data <= 8'b00000000 ;
			15'h00003A50 : data <= 8'b00000000 ;
			15'h00003A51 : data <= 8'b00000000 ;
			15'h00003A52 : data <= 8'b00000000 ;
			15'h00003A53 : data <= 8'b00000000 ;
			15'h00003A54 : data <= 8'b00000000 ;
			15'h00003A55 : data <= 8'b00000000 ;
			15'h00003A56 : data <= 8'b00000000 ;
			15'h00003A57 : data <= 8'b00000000 ;
			15'h00003A58 : data <= 8'b00000000 ;
			15'h00003A59 : data <= 8'b00000000 ;
			15'h00003A5A : data <= 8'b00000000 ;
			15'h00003A5B : data <= 8'b00000000 ;
			15'h00003A5C : data <= 8'b00000000 ;
			15'h00003A5D : data <= 8'b00000000 ;
			15'h00003A5E : data <= 8'b00000000 ;
			15'h00003A5F : data <= 8'b00000000 ;
			15'h00003A60 : data <= 8'b00000000 ;
			15'h00003A61 : data <= 8'b00000000 ;
			15'h00003A62 : data <= 8'b00000000 ;
			15'h00003A63 : data <= 8'b00000000 ;
			15'h00003A64 : data <= 8'b00000000 ;
			15'h00003A65 : data <= 8'b00000000 ;
			15'h00003A66 : data <= 8'b00000000 ;
			15'h00003A67 : data <= 8'b00000000 ;
			15'h00003A68 : data <= 8'b00000000 ;
			15'h00003A69 : data <= 8'b00000000 ;
			15'h00003A6A : data <= 8'b00000000 ;
			15'h00003A6B : data <= 8'b00000000 ;
			15'h00003A6C : data <= 8'b00000000 ;
			15'h00003A6D : data <= 8'b00000000 ;
			15'h00003A6E : data <= 8'b00000000 ;
			15'h00003A6F : data <= 8'b00000000 ;
			15'h00003A70 : data <= 8'b00000000 ;
			15'h00003A71 : data <= 8'b00000000 ;
			15'h00003A72 : data <= 8'b00000000 ;
			15'h00003A73 : data <= 8'b00000000 ;
			15'h00003A74 : data <= 8'b00000000 ;
			15'h00003A75 : data <= 8'b00000000 ;
			15'h00003A76 : data <= 8'b00000000 ;
			15'h00003A77 : data <= 8'b00000000 ;
			15'h00003A78 : data <= 8'b00000000 ;
			15'h00003A79 : data <= 8'b00000000 ;
			15'h00003A7A : data <= 8'b00000000 ;
			15'h00003A7B : data <= 8'b00000000 ;
			15'h00003A7C : data <= 8'b00000000 ;
			15'h00003A7D : data <= 8'b00000000 ;
			15'h00003A7E : data <= 8'b00000000 ;
			15'h00003A7F : data <= 8'b00000000 ;
			15'h00003A80 : data <= 8'b00000000 ;
			15'h00003A81 : data <= 8'b00000000 ;
			15'h00003A82 : data <= 8'b00000000 ;
			15'h00003A83 : data <= 8'b00000000 ;
			15'h00003A84 : data <= 8'b00000000 ;
			15'h00003A85 : data <= 8'b00000000 ;
			15'h00003A86 : data <= 8'b00000000 ;
			15'h00003A87 : data <= 8'b00000000 ;
			15'h00003A88 : data <= 8'b00000000 ;
			15'h00003A89 : data <= 8'b00000000 ;
			15'h00003A8A : data <= 8'b00000000 ;
			15'h00003A8B : data <= 8'b00000000 ;
			15'h00003A8C : data <= 8'b00000000 ;
			15'h00003A8D : data <= 8'b00000000 ;
			15'h00003A8E : data <= 8'b00000000 ;
			15'h00003A8F : data <= 8'b00000000 ;
			15'h00003A90 : data <= 8'b00000000 ;
			15'h00003A91 : data <= 8'b00000000 ;
			15'h00003A92 : data <= 8'b00000000 ;
			15'h00003A93 : data <= 8'b00000000 ;
			15'h00003A94 : data <= 8'b00000000 ;
			15'h00003A95 : data <= 8'b00000000 ;
			15'h00003A96 : data <= 8'b00000000 ;
			15'h00003A97 : data <= 8'b00000000 ;
			15'h00003A98 : data <= 8'b00000000 ;
			15'h00003A99 : data <= 8'b00000000 ;
			15'h00003A9A : data <= 8'b00000000 ;
			15'h00003A9B : data <= 8'b00000000 ;
			15'h00003A9C : data <= 8'b00000000 ;
			15'h00003A9D : data <= 8'b00000000 ;
			15'h00003A9E : data <= 8'b00000000 ;
			15'h00003A9F : data <= 8'b00000000 ;
			15'h00003AA0 : data <= 8'b00000000 ;
			15'h00003AA1 : data <= 8'b00000000 ;
			15'h00003AA2 : data <= 8'b00000000 ;
			15'h00003AA3 : data <= 8'b00000000 ;
			15'h00003AA4 : data <= 8'b00000000 ;
			15'h00003AA5 : data <= 8'b00000000 ;
			15'h00003AA6 : data <= 8'b00000000 ;
			15'h00003AA7 : data <= 8'b00000000 ;
			15'h00003AA8 : data <= 8'b00000000 ;
			15'h00003AA9 : data <= 8'b00000000 ;
			15'h00003AAA : data <= 8'b00000000 ;
			15'h00003AAB : data <= 8'b00000000 ;
			15'h00003AAC : data <= 8'b00000000 ;
			15'h00003AAD : data <= 8'b00000000 ;
			15'h00003AAE : data <= 8'b00000000 ;
			15'h00003AAF : data <= 8'b00000000 ;
			15'h00003AB0 : data <= 8'b00000000 ;
			15'h00003AB1 : data <= 8'b00000000 ;
			15'h00003AB2 : data <= 8'b00000000 ;
			15'h00003AB3 : data <= 8'b00000000 ;
			15'h00003AB4 : data <= 8'b00000000 ;
			15'h00003AB5 : data <= 8'b00000000 ;
			15'h00003AB6 : data <= 8'b00000000 ;
			15'h00003AB7 : data <= 8'b00000000 ;
			15'h00003AB8 : data <= 8'b00000000 ;
			15'h00003AB9 : data <= 8'b00000000 ;
			15'h00003ABA : data <= 8'b00000000 ;
			15'h00003ABB : data <= 8'b00000000 ;
			15'h00003ABC : data <= 8'b00000000 ;
			15'h00003ABD : data <= 8'b00000000 ;
			15'h00003ABE : data <= 8'b00000000 ;
			15'h00003ABF : data <= 8'b00000000 ;
			15'h00003AC0 : data <= 8'b00000000 ;
			15'h00003AC1 : data <= 8'b00000000 ;
			15'h00003AC2 : data <= 8'b00000000 ;
			15'h00003AC3 : data <= 8'b00000000 ;
			15'h00003AC4 : data <= 8'b00000000 ;
			15'h00003AC5 : data <= 8'b00000000 ;
			15'h00003AC6 : data <= 8'b00000000 ;
			15'h00003AC7 : data <= 8'b00000000 ;
			15'h00003AC8 : data <= 8'b00000000 ;
			15'h00003AC9 : data <= 8'b00000000 ;
			15'h00003ACA : data <= 8'b00000000 ;
			15'h00003ACB : data <= 8'b00000000 ;
			15'h00003ACC : data <= 8'b00000000 ;
			15'h00003ACD : data <= 8'b00000000 ;
			15'h00003ACE : data <= 8'b00000000 ;
			15'h00003ACF : data <= 8'b00000000 ;
			15'h00003AD0 : data <= 8'b00000000 ;
			15'h00003AD1 : data <= 8'b00000000 ;
			15'h00003AD2 : data <= 8'b00000000 ;
			15'h00003AD3 : data <= 8'b00000000 ;
			15'h00003AD4 : data <= 8'b00000000 ;
			15'h00003AD5 : data <= 8'b00000000 ;
			15'h00003AD6 : data <= 8'b00000000 ;
			15'h00003AD7 : data <= 8'b00000000 ;
			15'h00003AD8 : data <= 8'b00000000 ;
			15'h00003AD9 : data <= 8'b00000000 ;
			15'h00003ADA : data <= 8'b00000000 ;
			15'h00003ADB : data <= 8'b00000000 ;
			15'h00003ADC : data <= 8'b00000000 ;
			15'h00003ADD : data <= 8'b00000000 ;
			15'h00003ADE : data <= 8'b00000000 ;
			15'h00003ADF : data <= 8'b00000000 ;
			15'h00003AE0 : data <= 8'b00000000 ;
			15'h00003AE1 : data <= 8'b00000000 ;
			15'h00003AE2 : data <= 8'b00000000 ;
			15'h00003AE3 : data <= 8'b00000000 ;
			15'h00003AE4 : data <= 8'b00000000 ;
			15'h00003AE5 : data <= 8'b00000000 ;
			15'h00003AE6 : data <= 8'b00000000 ;
			15'h00003AE7 : data <= 8'b00000000 ;
			15'h00003AE8 : data <= 8'b00000000 ;
			15'h00003AE9 : data <= 8'b00000000 ;
			15'h00003AEA : data <= 8'b00000000 ;
			15'h00003AEB : data <= 8'b00000000 ;
			15'h00003AEC : data <= 8'b00000000 ;
			15'h00003AED : data <= 8'b00000000 ;
			15'h00003AEE : data <= 8'b00000000 ;
			15'h00003AEF : data <= 8'b00000000 ;
			15'h00003AF0 : data <= 8'b00000000 ;
			15'h00003AF1 : data <= 8'b00000000 ;
			15'h00003AF2 : data <= 8'b00000000 ;
			15'h00003AF3 : data <= 8'b00000000 ;
			15'h00003AF4 : data <= 8'b00000000 ;
			15'h00003AF5 : data <= 8'b00000000 ;
			15'h00003AF6 : data <= 8'b00000000 ;
			15'h00003AF7 : data <= 8'b00000000 ;
			15'h00003AF8 : data <= 8'b00000000 ;
			15'h00003AF9 : data <= 8'b00000000 ;
			15'h00003AFA : data <= 8'b00000000 ;
			15'h00003AFB : data <= 8'b00000000 ;
			15'h00003AFC : data <= 8'b00000000 ;
			15'h00003AFD : data <= 8'b00000000 ;
			15'h00003AFE : data <= 8'b00000000 ;
			15'h00003AFF : data <= 8'b00000000 ;
			15'h00003B00 : data <= 8'b00000000 ;
			15'h00003B01 : data <= 8'b00000000 ;
			15'h00003B02 : data <= 8'b00000000 ;
			15'h00003B03 : data <= 8'b00000000 ;
			15'h00003B04 : data <= 8'b00000000 ;
			15'h00003B05 : data <= 8'b00000000 ;
			15'h00003B06 : data <= 8'b00000000 ;
			15'h00003B07 : data <= 8'b00000000 ;
			15'h00003B08 : data <= 8'b00000000 ;
			15'h00003B09 : data <= 8'b00000000 ;
			15'h00003B0A : data <= 8'b00000000 ;
			15'h00003B0B : data <= 8'b00000000 ;
			15'h00003B0C : data <= 8'b00000000 ;
			15'h00003B0D : data <= 8'b00000000 ;
			15'h00003B0E : data <= 8'b00000000 ;
			15'h00003B0F : data <= 8'b00000000 ;
			15'h00003B10 : data <= 8'b00000000 ;
			15'h00003B11 : data <= 8'b00000000 ;
			15'h00003B12 : data <= 8'b00000000 ;
			15'h00003B13 : data <= 8'b00000000 ;
			15'h00003B14 : data <= 8'b00000000 ;
			15'h00003B15 : data <= 8'b00000000 ;
			15'h00003B16 : data <= 8'b00000000 ;
			15'h00003B17 : data <= 8'b00000000 ;
			15'h00003B18 : data <= 8'b00000000 ;
			15'h00003B19 : data <= 8'b00000000 ;
			15'h00003B1A : data <= 8'b00000000 ;
			15'h00003B1B : data <= 8'b00000000 ;
			15'h00003B1C : data <= 8'b00000000 ;
			15'h00003B1D : data <= 8'b00000000 ;
			15'h00003B1E : data <= 8'b00000000 ;
			15'h00003B1F : data <= 8'b00000000 ;
			15'h00003B20 : data <= 8'b00000000 ;
			15'h00003B21 : data <= 8'b00000000 ;
			15'h00003B22 : data <= 8'b00000000 ;
			15'h00003B23 : data <= 8'b00000000 ;
			15'h00003B24 : data <= 8'b00000000 ;
			15'h00003B25 : data <= 8'b00000000 ;
			15'h00003B26 : data <= 8'b00000000 ;
			15'h00003B27 : data <= 8'b00000000 ;
			15'h00003B28 : data <= 8'b00000000 ;
			15'h00003B29 : data <= 8'b00000000 ;
			15'h00003B2A : data <= 8'b00000000 ;
			15'h00003B2B : data <= 8'b00000000 ;
			15'h00003B2C : data <= 8'b00000000 ;
			15'h00003B2D : data <= 8'b00000000 ;
			15'h00003B2E : data <= 8'b00000000 ;
			15'h00003B2F : data <= 8'b00000000 ;
			15'h00003B30 : data <= 8'b00000000 ;
			15'h00003B31 : data <= 8'b00000000 ;
			15'h00003B32 : data <= 8'b00000000 ;
			15'h00003B33 : data <= 8'b00000000 ;
			15'h00003B34 : data <= 8'b00000000 ;
			15'h00003B35 : data <= 8'b00000000 ;
			15'h00003B36 : data <= 8'b00000000 ;
			15'h00003B37 : data <= 8'b00000000 ;
			15'h00003B38 : data <= 8'b00000000 ;
			15'h00003B39 : data <= 8'b00000000 ;
			15'h00003B3A : data <= 8'b00000000 ;
			15'h00003B3B : data <= 8'b00000000 ;
			15'h00003B3C : data <= 8'b00000000 ;
			15'h00003B3D : data <= 8'b00000000 ;
			15'h00003B3E : data <= 8'b00000000 ;
			15'h00003B3F : data <= 8'b00000000 ;
			15'h00003B40 : data <= 8'b00000000 ;
			15'h00003B41 : data <= 8'b00000000 ;
			15'h00003B42 : data <= 8'b00000000 ;
			15'h00003B43 : data <= 8'b00000000 ;
			15'h00003B44 : data <= 8'b00000000 ;
			15'h00003B45 : data <= 8'b00000000 ;
			15'h00003B46 : data <= 8'b00000000 ;
			15'h00003B47 : data <= 8'b00000000 ;
			15'h00003B48 : data <= 8'b00000000 ;
			15'h00003B49 : data <= 8'b00000000 ;
			15'h00003B4A : data <= 8'b00000000 ;
			15'h00003B4B : data <= 8'b00000000 ;
			15'h00003B4C : data <= 8'b00000000 ;
			15'h00003B4D : data <= 8'b00000000 ;
			15'h00003B4E : data <= 8'b00000000 ;
			15'h00003B4F : data <= 8'b00000000 ;
			15'h00003B50 : data <= 8'b00000000 ;
			15'h00003B51 : data <= 8'b00000000 ;
			15'h00003B52 : data <= 8'b00000000 ;
			15'h00003B53 : data <= 8'b00000000 ;
			15'h00003B54 : data <= 8'b00000000 ;
			15'h00003B55 : data <= 8'b00000000 ;
			15'h00003B56 : data <= 8'b00000000 ;
			15'h00003B57 : data <= 8'b00000000 ;
			15'h00003B58 : data <= 8'b00000000 ;
			15'h00003B59 : data <= 8'b00000000 ;
			15'h00003B5A : data <= 8'b00000000 ;
			15'h00003B5B : data <= 8'b00000000 ;
			15'h00003B5C : data <= 8'b00000000 ;
			15'h00003B5D : data <= 8'b00000000 ;
			15'h00003B5E : data <= 8'b00000000 ;
			15'h00003B5F : data <= 8'b00000000 ;
			15'h00003B60 : data <= 8'b00000000 ;
			15'h00003B61 : data <= 8'b00000000 ;
			15'h00003B62 : data <= 8'b00000000 ;
			15'h00003B63 : data <= 8'b00000000 ;
			15'h00003B64 : data <= 8'b00000000 ;
			15'h00003B65 : data <= 8'b00000000 ;
			15'h00003B66 : data <= 8'b00000000 ;
			15'h00003B67 : data <= 8'b00000000 ;
			15'h00003B68 : data <= 8'b00000000 ;
			15'h00003B69 : data <= 8'b00000000 ;
			15'h00003B6A : data <= 8'b00000000 ;
			15'h00003B6B : data <= 8'b00000000 ;
			15'h00003B6C : data <= 8'b00000000 ;
			15'h00003B6D : data <= 8'b00000000 ;
			15'h00003B6E : data <= 8'b00000000 ;
			15'h00003B6F : data <= 8'b00000000 ;
			15'h00003B70 : data <= 8'b00000000 ;
			15'h00003B71 : data <= 8'b00000000 ;
			15'h00003B72 : data <= 8'b00000000 ;
			15'h00003B73 : data <= 8'b00000000 ;
			15'h00003B74 : data <= 8'b00000000 ;
			15'h00003B75 : data <= 8'b00000000 ;
			15'h00003B76 : data <= 8'b00000000 ;
			15'h00003B77 : data <= 8'b00000000 ;
			15'h00003B78 : data <= 8'b00000000 ;
			15'h00003B79 : data <= 8'b00000000 ;
			15'h00003B7A : data <= 8'b00000000 ;
			15'h00003B7B : data <= 8'b00000000 ;
			15'h00003B7C : data <= 8'b00000000 ;
			15'h00003B7D : data <= 8'b00000000 ;
			15'h00003B7E : data <= 8'b00000000 ;
			15'h00003B7F : data <= 8'b00000000 ;
			15'h00003B80 : data <= 8'b00000000 ;
			15'h00003B81 : data <= 8'b00000000 ;
			15'h00003B82 : data <= 8'b00000000 ;
			15'h00003B83 : data <= 8'b00000000 ;
			15'h00003B84 : data <= 8'b00000000 ;
			15'h00003B85 : data <= 8'b00000000 ;
			15'h00003B86 : data <= 8'b00000000 ;
			15'h00003B87 : data <= 8'b00000000 ;
			15'h00003B88 : data <= 8'b00000000 ;
			15'h00003B89 : data <= 8'b00000000 ;
			15'h00003B8A : data <= 8'b00000000 ;
			15'h00003B8B : data <= 8'b00000000 ;
			15'h00003B8C : data <= 8'b00000000 ;
			15'h00003B8D : data <= 8'b00000000 ;
			15'h00003B8E : data <= 8'b00000000 ;
			15'h00003B8F : data <= 8'b00000000 ;
			15'h00003B90 : data <= 8'b00000000 ;
			15'h00003B91 : data <= 8'b00000000 ;
			15'h00003B92 : data <= 8'b00000000 ;
			15'h00003B93 : data <= 8'b00000000 ;
			15'h00003B94 : data <= 8'b00000000 ;
			15'h00003B95 : data <= 8'b00000000 ;
			15'h00003B96 : data <= 8'b00000000 ;
			15'h00003B97 : data <= 8'b00000000 ;
			15'h00003B98 : data <= 8'b00000000 ;
			15'h00003B99 : data <= 8'b00000000 ;
			15'h00003B9A : data <= 8'b00000000 ;
			15'h00003B9B : data <= 8'b00000000 ;
			15'h00003B9C : data <= 8'b00000000 ;
			15'h00003B9D : data <= 8'b00000000 ;
			15'h00003B9E : data <= 8'b00000000 ;
			15'h00003B9F : data <= 8'b00000000 ;
			15'h00003BA0 : data <= 8'b00000000 ;
			15'h00003BA1 : data <= 8'b00000000 ;
			15'h00003BA2 : data <= 8'b00000000 ;
			15'h00003BA3 : data <= 8'b00000000 ;
			15'h00003BA4 : data <= 8'b00000000 ;
			15'h00003BA5 : data <= 8'b00000000 ;
			15'h00003BA6 : data <= 8'b00000000 ;
			15'h00003BA7 : data <= 8'b00000000 ;
			15'h00003BA8 : data <= 8'b00000000 ;
			15'h00003BA9 : data <= 8'b00000000 ;
			15'h00003BAA : data <= 8'b00000000 ;
			15'h00003BAB : data <= 8'b00000000 ;
			15'h00003BAC : data <= 8'b00000000 ;
			15'h00003BAD : data <= 8'b00000000 ;
			15'h00003BAE : data <= 8'b00000000 ;
			15'h00003BAF : data <= 8'b00000000 ;
			15'h00003BB0 : data <= 8'b00000000 ;
			15'h00003BB1 : data <= 8'b00000000 ;
			15'h00003BB2 : data <= 8'b00000000 ;
			15'h00003BB3 : data <= 8'b00000000 ;
			15'h00003BB4 : data <= 8'b00000000 ;
			15'h00003BB5 : data <= 8'b00000000 ;
			15'h00003BB6 : data <= 8'b00000000 ;
			15'h00003BB7 : data <= 8'b00000000 ;
			15'h00003BB8 : data <= 8'b00000000 ;
			15'h00003BB9 : data <= 8'b00000000 ;
			15'h00003BBA : data <= 8'b00000000 ;
			15'h00003BBB : data <= 8'b00000000 ;
			15'h00003BBC : data <= 8'b00000000 ;
			15'h00003BBD : data <= 8'b00000000 ;
			15'h00003BBE : data <= 8'b00000000 ;
			15'h00003BBF : data <= 8'b00000000 ;
			15'h00003BC0 : data <= 8'b00000000 ;
			15'h00003BC1 : data <= 8'b00000000 ;
			15'h00003BC2 : data <= 8'b00000000 ;
			15'h00003BC3 : data <= 8'b00000000 ;
			15'h00003BC4 : data <= 8'b00000000 ;
			15'h00003BC5 : data <= 8'b00000000 ;
			15'h00003BC6 : data <= 8'b00000000 ;
			15'h00003BC7 : data <= 8'b00000000 ;
			15'h00003BC8 : data <= 8'b00000000 ;
			15'h00003BC9 : data <= 8'b00000000 ;
			15'h00003BCA : data <= 8'b00000000 ;
			15'h00003BCB : data <= 8'b00000000 ;
			15'h00003BCC : data <= 8'b00000000 ;
			15'h00003BCD : data <= 8'b00000000 ;
			15'h00003BCE : data <= 8'b00000000 ;
			15'h00003BCF : data <= 8'b00000000 ;
			15'h00003BD0 : data <= 8'b00000000 ;
			15'h00003BD1 : data <= 8'b00000000 ;
			15'h00003BD2 : data <= 8'b00000000 ;
			15'h00003BD3 : data <= 8'b00000000 ;
			15'h00003BD4 : data <= 8'b00000000 ;
			15'h00003BD5 : data <= 8'b00000000 ;
			15'h00003BD6 : data <= 8'b00000000 ;
			15'h00003BD7 : data <= 8'b00000000 ;
			15'h00003BD8 : data <= 8'b00000000 ;
			15'h00003BD9 : data <= 8'b00000000 ;
			15'h00003BDA : data <= 8'b00000000 ;
			15'h00003BDB : data <= 8'b00000000 ;
			15'h00003BDC : data <= 8'b00000000 ;
			15'h00003BDD : data <= 8'b00000000 ;
			15'h00003BDE : data <= 8'b00000000 ;
			15'h00003BDF : data <= 8'b00000000 ;
			15'h00003BE0 : data <= 8'b00000000 ;
			15'h00003BE1 : data <= 8'b00000000 ;
			15'h00003BE2 : data <= 8'b00000000 ;
			15'h00003BE3 : data <= 8'b00000000 ;
			15'h00003BE4 : data <= 8'b00000000 ;
			15'h00003BE5 : data <= 8'b00000000 ;
			15'h00003BE6 : data <= 8'b00000000 ;
			15'h00003BE7 : data <= 8'b00000000 ;
			15'h00003BE8 : data <= 8'b00000000 ;
			15'h00003BE9 : data <= 8'b00000000 ;
			15'h00003BEA : data <= 8'b00000000 ;
			15'h00003BEB : data <= 8'b00000000 ;
			15'h00003BEC : data <= 8'b00000000 ;
			15'h00003BED : data <= 8'b00000000 ;
			15'h00003BEE : data <= 8'b00000000 ;
			15'h00003BEF : data <= 8'b00000000 ;
			15'h00003BF0 : data <= 8'b00000000 ;
			15'h00003BF1 : data <= 8'b00000000 ;
			15'h00003BF2 : data <= 8'b00000000 ;
			15'h00003BF3 : data <= 8'b00000000 ;
			15'h00003BF4 : data <= 8'b00000000 ;
			15'h00003BF5 : data <= 8'b00000000 ;
			15'h00003BF6 : data <= 8'b00000000 ;
			15'h00003BF7 : data <= 8'b00000000 ;
			15'h00003BF8 : data <= 8'b00000000 ;
			15'h00003BF9 : data <= 8'b00000000 ;
			15'h00003BFA : data <= 8'b00000000 ;
			15'h00003BFB : data <= 8'b00000000 ;
			15'h00003BFC : data <= 8'b00000000 ;
			15'h00003BFD : data <= 8'b00000000 ;
			15'h00003BFE : data <= 8'b00000000 ;
			15'h00003BFF : data <= 8'b00000000 ;
			15'h00003C00 : data <= 8'b00000000 ;
			15'h00003C01 : data <= 8'b00000000 ;
			15'h00003C02 : data <= 8'b00000000 ;
			15'h00003C03 : data <= 8'b00000000 ;
			15'h00003C04 : data <= 8'b00000000 ;
			15'h00003C05 : data <= 8'b00000000 ;
			15'h00003C06 : data <= 8'b00000000 ;
			15'h00003C07 : data <= 8'b00000000 ;
			15'h00003C08 : data <= 8'b00000000 ;
			15'h00003C09 : data <= 8'b00000000 ;
			15'h00003C0A : data <= 8'b00000000 ;
			15'h00003C0B : data <= 8'b00000000 ;
			15'h00003C0C : data <= 8'b00000000 ;
			15'h00003C0D : data <= 8'b00000000 ;
			15'h00003C0E : data <= 8'b00000000 ;
			15'h00003C0F : data <= 8'b00000000 ;
			15'h00003C10 : data <= 8'b00000000 ;
			15'h00003C11 : data <= 8'b00000000 ;
			15'h00003C12 : data <= 8'b00000000 ;
			15'h00003C13 : data <= 8'b00000000 ;
			15'h00003C14 : data <= 8'b00000000 ;
			15'h00003C15 : data <= 8'b00000000 ;
			15'h00003C16 : data <= 8'b00000000 ;
			15'h00003C17 : data <= 8'b00000000 ;
			15'h00003C18 : data <= 8'b00000000 ;
			15'h00003C19 : data <= 8'b00000000 ;
			15'h00003C1A : data <= 8'b00000000 ;
			15'h00003C1B : data <= 8'b00000000 ;
			15'h00003C1C : data <= 8'b00000000 ;
			15'h00003C1D : data <= 8'b00000000 ;
			15'h00003C1E : data <= 8'b00000000 ;
			15'h00003C1F : data <= 8'b00000000 ;
			15'h00003C20 : data <= 8'b00000000 ;
			15'h00003C21 : data <= 8'b00000000 ;
			15'h00003C22 : data <= 8'b00000000 ;
			15'h00003C23 : data <= 8'b00000000 ;
			15'h00003C24 : data <= 8'b00000000 ;
			15'h00003C25 : data <= 8'b00000000 ;
			15'h00003C26 : data <= 8'b00000000 ;
			15'h00003C27 : data <= 8'b00000000 ;
			15'h00003C28 : data <= 8'b00000000 ;
			15'h00003C29 : data <= 8'b00000000 ;
			15'h00003C2A : data <= 8'b00000000 ;
			15'h00003C2B : data <= 8'b00000000 ;
			15'h00003C2C : data <= 8'b00000000 ;
			15'h00003C2D : data <= 8'b00000000 ;
			15'h00003C2E : data <= 8'b00000000 ;
			15'h00003C2F : data <= 8'b00000000 ;
			15'h00003C30 : data <= 8'b00000000 ;
			15'h00003C31 : data <= 8'b00000000 ;
			15'h00003C32 : data <= 8'b00000000 ;
			15'h00003C33 : data <= 8'b00000000 ;
			15'h00003C34 : data <= 8'b00000000 ;
			15'h00003C35 : data <= 8'b00000000 ;
			15'h00003C36 : data <= 8'b00000000 ;
			15'h00003C37 : data <= 8'b00000000 ;
			15'h00003C38 : data <= 8'b00000000 ;
			15'h00003C39 : data <= 8'b00000000 ;
			15'h00003C3A : data <= 8'b00000000 ;
			15'h00003C3B : data <= 8'b00000000 ;
			15'h00003C3C : data <= 8'b00000000 ;
			15'h00003C3D : data <= 8'b00000000 ;
			15'h00003C3E : data <= 8'b00000000 ;
			15'h00003C3F : data <= 8'b00000000 ;
			15'h00003C40 : data <= 8'b00000000 ;
			15'h00003C41 : data <= 8'b00000000 ;
			15'h00003C42 : data <= 8'b00000000 ;
			15'h00003C43 : data <= 8'b00000000 ;
			15'h00003C44 : data <= 8'b00000000 ;
			15'h00003C45 : data <= 8'b00000000 ;
			15'h00003C46 : data <= 8'b00000000 ;
			15'h00003C47 : data <= 8'b00000000 ;
			15'h00003C48 : data <= 8'b00000000 ;
			15'h00003C49 : data <= 8'b00000000 ;
			15'h00003C4A : data <= 8'b00000000 ;
			15'h00003C4B : data <= 8'b00000000 ;
			15'h00003C4C : data <= 8'b00000000 ;
			15'h00003C4D : data <= 8'b00000000 ;
			15'h00003C4E : data <= 8'b00000000 ;
			15'h00003C4F : data <= 8'b00000000 ;
			15'h00003C50 : data <= 8'b00000000 ;
			15'h00003C51 : data <= 8'b00000000 ;
			15'h00003C52 : data <= 8'b00000000 ;
			15'h00003C53 : data <= 8'b00000000 ;
			15'h00003C54 : data <= 8'b00000000 ;
			15'h00003C55 : data <= 8'b00000000 ;
			15'h00003C56 : data <= 8'b00000000 ;
			15'h00003C57 : data <= 8'b00000000 ;
			15'h00003C58 : data <= 8'b00000000 ;
			15'h00003C59 : data <= 8'b00000000 ;
			15'h00003C5A : data <= 8'b00000000 ;
			15'h00003C5B : data <= 8'b00000000 ;
			15'h00003C5C : data <= 8'b00000000 ;
			15'h00003C5D : data <= 8'b00000000 ;
			15'h00003C5E : data <= 8'b00000000 ;
			15'h00003C5F : data <= 8'b00000000 ;
			15'h00003C60 : data <= 8'b00000000 ;
			15'h00003C61 : data <= 8'b00000000 ;
			15'h00003C62 : data <= 8'b00000000 ;
			15'h00003C63 : data <= 8'b00000000 ;
			15'h00003C64 : data <= 8'b00000000 ;
			15'h00003C65 : data <= 8'b00000000 ;
			15'h00003C66 : data <= 8'b00000000 ;
			15'h00003C67 : data <= 8'b00000000 ;
			15'h00003C68 : data <= 8'b00000000 ;
			15'h00003C69 : data <= 8'b00000000 ;
			15'h00003C6A : data <= 8'b00000000 ;
			15'h00003C6B : data <= 8'b00000000 ;
			15'h00003C6C : data <= 8'b00000000 ;
			15'h00003C6D : data <= 8'b00000000 ;
			15'h00003C6E : data <= 8'b00000000 ;
			15'h00003C6F : data <= 8'b00000000 ;
			15'h00003C70 : data <= 8'b00000000 ;
			15'h00003C71 : data <= 8'b00000000 ;
			15'h00003C72 : data <= 8'b00000000 ;
			15'h00003C73 : data <= 8'b00000000 ;
			15'h00003C74 : data <= 8'b00000000 ;
			15'h00003C75 : data <= 8'b00000000 ;
			15'h00003C76 : data <= 8'b00000000 ;
			15'h00003C77 : data <= 8'b00000000 ;
			15'h00003C78 : data <= 8'b00000000 ;
			15'h00003C79 : data <= 8'b00000000 ;
			15'h00003C7A : data <= 8'b00000000 ;
			15'h00003C7B : data <= 8'b00000000 ;
			15'h00003C7C : data <= 8'b00000000 ;
			15'h00003C7D : data <= 8'b00000000 ;
			15'h00003C7E : data <= 8'b00000000 ;
			15'h00003C7F : data <= 8'b00000000 ;
			15'h00003C80 : data <= 8'b00000000 ;
			15'h00003C81 : data <= 8'b00000000 ;
			15'h00003C82 : data <= 8'b00000000 ;
			15'h00003C83 : data <= 8'b00000000 ;
			15'h00003C84 : data <= 8'b00000000 ;
			15'h00003C85 : data <= 8'b00000000 ;
			15'h00003C86 : data <= 8'b00000000 ;
			15'h00003C87 : data <= 8'b00000000 ;
			15'h00003C88 : data <= 8'b00000000 ;
			15'h00003C89 : data <= 8'b00000000 ;
			15'h00003C8A : data <= 8'b00000000 ;
			15'h00003C8B : data <= 8'b00000000 ;
			15'h00003C8C : data <= 8'b00000000 ;
			15'h00003C8D : data <= 8'b00000000 ;
			15'h00003C8E : data <= 8'b00000000 ;
			15'h00003C8F : data <= 8'b00000000 ;
			15'h00003C90 : data <= 8'b00000000 ;
			15'h00003C91 : data <= 8'b00000000 ;
			15'h00003C92 : data <= 8'b00000000 ;
			15'h00003C93 : data <= 8'b00000000 ;
			15'h00003C94 : data <= 8'b00000000 ;
			15'h00003C95 : data <= 8'b00000000 ;
			15'h00003C96 : data <= 8'b00000000 ;
			15'h00003C97 : data <= 8'b00000000 ;
			15'h00003C98 : data <= 8'b00000000 ;
			15'h00003C99 : data <= 8'b00000000 ;
			15'h00003C9A : data <= 8'b00000000 ;
			15'h00003C9B : data <= 8'b00000000 ;
			15'h00003C9C : data <= 8'b00000000 ;
			15'h00003C9D : data <= 8'b00000000 ;
			15'h00003C9E : data <= 8'b00000000 ;
			15'h00003C9F : data <= 8'b00000000 ;
			15'h00003CA0 : data <= 8'b00000000 ;
			15'h00003CA1 : data <= 8'b00000000 ;
			15'h00003CA2 : data <= 8'b00000000 ;
			15'h00003CA3 : data <= 8'b00000000 ;
			15'h00003CA4 : data <= 8'b00000000 ;
			15'h00003CA5 : data <= 8'b00000000 ;
			15'h00003CA6 : data <= 8'b00000000 ;
			15'h00003CA7 : data <= 8'b00000000 ;
			15'h00003CA8 : data <= 8'b00000000 ;
			15'h00003CA9 : data <= 8'b00000000 ;
			15'h00003CAA : data <= 8'b00000000 ;
			15'h00003CAB : data <= 8'b00000000 ;
			15'h00003CAC : data <= 8'b00000000 ;
			15'h00003CAD : data <= 8'b00000000 ;
			15'h00003CAE : data <= 8'b00000000 ;
			15'h00003CAF : data <= 8'b00000000 ;
			15'h00003CB0 : data <= 8'b00000000 ;
			15'h00003CB1 : data <= 8'b00000000 ;
			15'h00003CB2 : data <= 8'b00000000 ;
			15'h00003CB3 : data <= 8'b00000000 ;
			15'h00003CB4 : data <= 8'b00000000 ;
			15'h00003CB5 : data <= 8'b00000000 ;
			15'h00003CB6 : data <= 8'b00000000 ;
			15'h00003CB7 : data <= 8'b00000000 ;
			15'h00003CB8 : data <= 8'b00000000 ;
			15'h00003CB9 : data <= 8'b00000000 ;
			15'h00003CBA : data <= 8'b00000000 ;
			15'h00003CBB : data <= 8'b00000000 ;
			15'h00003CBC : data <= 8'b00000000 ;
			15'h00003CBD : data <= 8'b00000000 ;
			15'h00003CBE : data <= 8'b00000000 ;
			15'h00003CBF : data <= 8'b00000000 ;
			15'h00003CC0 : data <= 8'b00000000 ;
			15'h00003CC1 : data <= 8'b00000000 ;
			15'h00003CC2 : data <= 8'b00000000 ;
			15'h00003CC3 : data <= 8'b00000000 ;
			15'h00003CC4 : data <= 8'b00000000 ;
			15'h00003CC5 : data <= 8'b00000000 ;
			15'h00003CC6 : data <= 8'b00000000 ;
			15'h00003CC7 : data <= 8'b00000000 ;
			15'h00003CC8 : data <= 8'b00000000 ;
			15'h00003CC9 : data <= 8'b00000000 ;
			15'h00003CCA : data <= 8'b00000000 ;
			15'h00003CCB : data <= 8'b00000000 ;
			15'h00003CCC : data <= 8'b00000000 ;
			15'h00003CCD : data <= 8'b00000000 ;
			15'h00003CCE : data <= 8'b00000000 ;
			15'h00003CCF : data <= 8'b00000000 ;
			15'h00003CD0 : data <= 8'b00000000 ;
			15'h00003CD1 : data <= 8'b00000000 ;
			15'h00003CD2 : data <= 8'b00000000 ;
			15'h00003CD3 : data <= 8'b00000000 ;
			15'h00003CD4 : data <= 8'b00000000 ;
			15'h00003CD5 : data <= 8'b00000000 ;
			15'h00003CD6 : data <= 8'b00000000 ;
			15'h00003CD7 : data <= 8'b00000000 ;
			15'h00003CD8 : data <= 8'b00000000 ;
			15'h00003CD9 : data <= 8'b00000000 ;
			15'h00003CDA : data <= 8'b00000000 ;
			15'h00003CDB : data <= 8'b00000000 ;
			15'h00003CDC : data <= 8'b00000000 ;
			15'h00003CDD : data <= 8'b00000000 ;
			15'h00003CDE : data <= 8'b00000000 ;
			15'h00003CDF : data <= 8'b00000000 ;
			15'h00003CE0 : data <= 8'b00000000 ;
			15'h00003CE1 : data <= 8'b00000000 ;
			15'h00003CE2 : data <= 8'b00000000 ;
			15'h00003CE3 : data <= 8'b00000000 ;
			15'h00003CE4 : data <= 8'b00000000 ;
			15'h00003CE5 : data <= 8'b00000000 ;
			15'h00003CE6 : data <= 8'b00000000 ;
			15'h00003CE7 : data <= 8'b00000000 ;
			15'h00003CE8 : data <= 8'b00000000 ;
			15'h00003CE9 : data <= 8'b00000000 ;
			15'h00003CEA : data <= 8'b00000000 ;
			15'h00003CEB : data <= 8'b00000000 ;
			15'h00003CEC : data <= 8'b00000000 ;
			15'h00003CED : data <= 8'b00000000 ;
			15'h00003CEE : data <= 8'b00000000 ;
			15'h00003CEF : data <= 8'b00000000 ;
			15'h00003CF0 : data <= 8'b00000000 ;
			15'h00003CF1 : data <= 8'b00000000 ;
			15'h00003CF2 : data <= 8'b00000000 ;
			15'h00003CF3 : data <= 8'b00000000 ;
			15'h00003CF4 : data <= 8'b00000000 ;
			15'h00003CF5 : data <= 8'b00000000 ;
			15'h00003CF6 : data <= 8'b00000000 ;
			15'h00003CF7 : data <= 8'b00000000 ;
			15'h00003CF8 : data <= 8'b00000000 ;
			15'h00003CF9 : data <= 8'b00000000 ;
			15'h00003CFA : data <= 8'b00000000 ;
			15'h00003CFB : data <= 8'b00000000 ;
			15'h00003CFC : data <= 8'b00000000 ;
			15'h00003CFD : data <= 8'b00000000 ;
			15'h00003CFE : data <= 8'b00000000 ;
			15'h00003CFF : data <= 8'b00000000 ;
			15'h00003D00 : data <= 8'b00000000 ;
			15'h00003D01 : data <= 8'b00000000 ;
			15'h00003D02 : data <= 8'b00000000 ;
			15'h00003D03 : data <= 8'b00000000 ;
			15'h00003D04 : data <= 8'b00000000 ;
			15'h00003D05 : data <= 8'b00000000 ;
			15'h00003D06 : data <= 8'b00000000 ;
			15'h00003D07 : data <= 8'b00000000 ;
			15'h00003D08 : data <= 8'b00000000 ;
			15'h00003D09 : data <= 8'b00000000 ;
			15'h00003D0A : data <= 8'b00000000 ;
			15'h00003D0B : data <= 8'b00000000 ;
			15'h00003D0C : data <= 8'b00000000 ;
			15'h00003D0D : data <= 8'b00000000 ;
			15'h00003D0E : data <= 8'b00000000 ;
			15'h00003D0F : data <= 8'b00000000 ;
			15'h00003D10 : data <= 8'b00000000 ;
			15'h00003D11 : data <= 8'b00000000 ;
			15'h00003D12 : data <= 8'b00000000 ;
			15'h00003D13 : data <= 8'b00000000 ;
			15'h00003D14 : data <= 8'b00000000 ;
			15'h00003D15 : data <= 8'b00000000 ;
			15'h00003D16 : data <= 8'b00000000 ;
			15'h00003D17 : data <= 8'b00000000 ;
			15'h00003D18 : data <= 8'b00000000 ;
			15'h00003D19 : data <= 8'b00000000 ;
			15'h00003D1A : data <= 8'b00000000 ;
			15'h00003D1B : data <= 8'b00000000 ;
			15'h00003D1C : data <= 8'b00000000 ;
			15'h00003D1D : data <= 8'b00000000 ;
			15'h00003D1E : data <= 8'b00000000 ;
			15'h00003D1F : data <= 8'b00000000 ;
			15'h00003D20 : data <= 8'b00000000 ;
			15'h00003D21 : data <= 8'b00000000 ;
			15'h00003D22 : data <= 8'b00000000 ;
			15'h00003D23 : data <= 8'b00000000 ;
			15'h00003D24 : data <= 8'b00000000 ;
			15'h00003D25 : data <= 8'b00000000 ;
			15'h00003D26 : data <= 8'b00000000 ;
			15'h00003D27 : data <= 8'b00000000 ;
			15'h00003D28 : data <= 8'b00000000 ;
			15'h00003D29 : data <= 8'b00000000 ;
			15'h00003D2A : data <= 8'b00000000 ;
			15'h00003D2B : data <= 8'b00000000 ;
			15'h00003D2C : data <= 8'b00000000 ;
			15'h00003D2D : data <= 8'b00000000 ;
			15'h00003D2E : data <= 8'b00000000 ;
			15'h00003D2F : data <= 8'b00000000 ;
			15'h00003D30 : data <= 8'b00000000 ;
			15'h00003D31 : data <= 8'b00000000 ;
			15'h00003D32 : data <= 8'b00000000 ;
			15'h00003D33 : data <= 8'b00000000 ;
			15'h00003D34 : data <= 8'b00000000 ;
			15'h00003D35 : data <= 8'b00000000 ;
			15'h00003D36 : data <= 8'b00000000 ;
			15'h00003D37 : data <= 8'b00000000 ;
			15'h00003D38 : data <= 8'b00000000 ;
			15'h00003D39 : data <= 8'b00000000 ;
			15'h00003D3A : data <= 8'b00000000 ;
			15'h00003D3B : data <= 8'b00000000 ;
			15'h00003D3C : data <= 8'b00000000 ;
			15'h00003D3D : data <= 8'b00000000 ;
			15'h00003D3E : data <= 8'b00000000 ;
			15'h00003D3F : data <= 8'b00000000 ;
			15'h00003D40 : data <= 8'b00000000 ;
			15'h00003D41 : data <= 8'b00000000 ;
			15'h00003D42 : data <= 8'b00000000 ;
			15'h00003D43 : data <= 8'b00000000 ;
			15'h00003D44 : data <= 8'b00000000 ;
			15'h00003D45 : data <= 8'b00000000 ;
			15'h00003D46 : data <= 8'b00000000 ;
			15'h00003D47 : data <= 8'b00000000 ;
			15'h00003D48 : data <= 8'b00000000 ;
			15'h00003D49 : data <= 8'b00000000 ;
			15'h00003D4A : data <= 8'b00000000 ;
			15'h00003D4B : data <= 8'b00000000 ;
			15'h00003D4C : data <= 8'b00000000 ;
			15'h00003D4D : data <= 8'b00000000 ;
			15'h00003D4E : data <= 8'b00000000 ;
			15'h00003D4F : data <= 8'b00000000 ;
			15'h00003D50 : data <= 8'b00000000 ;
			15'h00003D51 : data <= 8'b00000000 ;
			15'h00003D52 : data <= 8'b00000000 ;
			15'h00003D53 : data <= 8'b00000000 ;
			15'h00003D54 : data <= 8'b00000000 ;
			15'h00003D55 : data <= 8'b00000000 ;
			15'h00003D56 : data <= 8'b00000000 ;
			15'h00003D57 : data <= 8'b00000000 ;
			15'h00003D58 : data <= 8'b00000000 ;
			15'h00003D59 : data <= 8'b00000000 ;
			15'h00003D5A : data <= 8'b00000000 ;
			15'h00003D5B : data <= 8'b00000000 ;
			15'h00003D5C : data <= 8'b00000000 ;
			15'h00003D5D : data <= 8'b00000000 ;
			15'h00003D5E : data <= 8'b00000000 ;
			15'h00003D5F : data <= 8'b00000000 ;
			15'h00003D60 : data <= 8'b00000000 ;
			15'h00003D61 : data <= 8'b00000000 ;
			15'h00003D62 : data <= 8'b00000000 ;
			15'h00003D63 : data <= 8'b00000000 ;
			15'h00003D64 : data <= 8'b00000000 ;
			15'h00003D65 : data <= 8'b00000000 ;
			15'h00003D66 : data <= 8'b00000000 ;
			15'h00003D67 : data <= 8'b00000000 ;
			15'h00003D68 : data <= 8'b00000000 ;
			15'h00003D69 : data <= 8'b00000000 ;
			15'h00003D6A : data <= 8'b00000000 ;
			15'h00003D6B : data <= 8'b00000000 ;
			15'h00003D6C : data <= 8'b00000000 ;
			15'h00003D6D : data <= 8'b00000000 ;
			15'h00003D6E : data <= 8'b00000000 ;
			15'h00003D6F : data <= 8'b00000000 ;
			15'h00003D70 : data <= 8'b00000000 ;
			15'h00003D71 : data <= 8'b00000000 ;
			15'h00003D72 : data <= 8'b00000000 ;
			15'h00003D73 : data <= 8'b00000000 ;
			15'h00003D74 : data <= 8'b00000000 ;
			15'h00003D75 : data <= 8'b00000000 ;
			15'h00003D76 : data <= 8'b00000000 ;
			15'h00003D77 : data <= 8'b00000000 ;
			15'h00003D78 : data <= 8'b00000000 ;
			15'h00003D79 : data <= 8'b00000000 ;
			15'h00003D7A : data <= 8'b00000000 ;
			15'h00003D7B : data <= 8'b00000000 ;
			15'h00003D7C : data <= 8'b00000000 ;
			15'h00003D7D : data <= 8'b00000000 ;
			15'h00003D7E : data <= 8'b00000000 ;
			15'h00003D7F : data <= 8'b00000000 ;
			15'h00003D80 : data <= 8'b00000000 ;
			15'h00003D81 : data <= 8'b00000000 ;
			15'h00003D82 : data <= 8'b00000000 ;
			15'h00003D83 : data <= 8'b00000000 ;
			15'h00003D84 : data <= 8'b00000000 ;
			15'h00003D85 : data <= 8'b00000000 ;
			15'h00003D86 : data <= 8'b00000000 ;
			15'h00003D87 : data <= 8'b00000000 ;
			15'h00003D88 : data <= 8'b00000000 ;
			15'h00003D89 : data <= 8'b00000000 ;
			15'h00003D8A : data <= 8'b00000000 ;
			15'h00003D8B : data <= 8'b00000000 ;
			15'h00003D8C : data <= 8'b00000000 ;
			15'h00003D8D : data <= 8'b00000000 ;
			15'h00003D8E : data <= 8'b00000000 ;
			15'h00003D8F : data <= 8'b00000000 ;
			15'h00003D90 : data <= 8'b00000000 ;
			15'h00003D91 : data <= 8'b00000000 ;
			15'h00003D92 : data <= 8'b00000000 ;
			15'h00003D93 : data <= 8'b00000000 ;
			15'h00003D94 : data <= 8'b00000000 ;
			15'h00003D95 : data <= 8'b00000000 ;
			15'h00003D96 : data <= 8'b00000000 ;
			15'h00003D97 : data <= 8'b00000000 ;
			15'h00003D98 : data <= 8'b00000000 ;
			15'h00003D99 : data <= 8'b00000000 ;
			15'h00003D9A : data <= 8'b00000000 ;
			15'h00003D9B : data <= 8'b00000000 ;
			15'h00003D9C : data <= 8'b00000000 ;
			15'h00003D9D : data <= 8'b00000000 ;
			15'h00003D9E : data <= 8'b00000000 ;
			15'h00003D9F : data <= 8'b00000000 ;
			15'h00003DA0 : data <= 8'b00000000 ;
			15'h00003DA1 : data <= 8'b00000000 ;
			15'h00003DA2 : data <= 8'b00000000 ;
			15'h00003DA3 : data <= 8'b00000000 ;
			15'h00003DA4 : data <= 8'b00000000 ;
			15'h00003DA5 : data <= 8'b00000000 ;
			15'h00003DA6 : data <= 8'b00000000 ;
			15'h00003DA7 : data <= 8'b00000000 ;
			15'h00003DA8 : data <= 8'b00000000 ;
			15'h00003DA9 : data <= 8'b00000000 ;
			15'h00003DAA : data <= 8'b00000000 ;
			15'h00003DAB : data <= 8'b00000000 ;
			15'h00003DAC : data <= 8'b00000000 ;
			15'h00003DAD : data <= 8'b00000000 ;
			15'h00003DAE : data <= 8'b00000000 ;
			15'h00003DAF : data <= 8'b00000000 ;
			15'h00003DB0 : data <= 8'b00000000 ;
			15'h00003DB1 : data <= 8'b00000000 ;
			15'h00003DB2 : data <= 8'b00000000 ;
			15'h00003DB3 : data <= 8'b00000000 ;
			15'h00003DB4 : data <= 8'b00000000 ;
			15'h00003DB5 : data <= 8'b00000000 ;
			15'h00003DB6 : data <= 8'b00000000 ;
			15'h00003DB7 : data <= 8'b00000000 ;
			15'h00003DB8 : data <= 8'b00000000 ;
			15'h00003DB9 : data <= 8'b00000000 ;
			15'h00003DBA : data <= 8'b00000000 ;
			15'h00003DBB : data <= 8'b00000000 ;
			15'h00003DBC : data <= 8'b00000000 ;
			15'h00003DBD : data <= 8'b00000000 ;
			15'h00003DBE : data <= 8'b00000000 ;
			15'h00003DBF : data <= 8'b00000000 ;
			15'h00003DC0 : data <= 8'b00000000 ;
			15'h00003DC1 : data <= 8'b00000000 ;
			15'h00003DC2 : data <= 8'b00000000 ;
			15'h00003DC3 : data <= 8'b00000000 ;
			15'h00003DC4 : data <= 8'b00000000 ;
			15'h00003DC5 : data <= 8'b00000000 ;
			15'h00003DC6 : data <= 8'b00000000 ;
			15'h00003DC7 : data <= 8'b00000000 ;
			15'h00003DC8 : data <= 8'b00000000 ;
			15'h00003DC9 : data <= 8'b00000000 ;
			15'h00003DCA : data <= 8'b00000000 ;
			15'h00003DCB : data <= 8'b00000000 ;
			15'h00003DCC : data <= 8'b00000000 ;
			15'h00003DCD : data <= 8'b00000000 ;
			15'h00003DCE : data <= 8'b00000000 ;
			15'h00003DCF : data <= 8'b00000000 ;
			15'h00003DD0 : data <= 8'b00000000 ;
			15'h00003DD1 : data <= 8'b00000000 ;
			15'h00003DD2 : data <= 8'b00000000 ;
			15'h00003DD3 : data <= 8'b00000000 ;
			15'h00003DD4 : data <= 8'b00000000 ;
			15'h00003DD5 : data <= 8'b00000000 ;
			15'h00003DD6 : data <= 8'b00000000 ;
			15'h00003DD7 : data <= 8'b00000000 ;
			15'h00003DD8 : data <= 8'b00000000 ;
			15'h00003DD9 : data <= 8'b00000000 ;
			15'h00003DDA : data <= 8'b00000000 ;
			15'h00003DDB : data <= 8'b00000000 ;
			15'h00003DDC : data <= 8'b00000000 ;
			15'h00003DDD : data <= 8'b00000000 ;
			15'h00003DDE : data <= 8'b00000000 ;
			15'h00003DDF : data <= 8'b00000000 ;
			15'h00003DE0 : data <= 8'b00000000 ;
			15'h00003DE1 : data <= 8'b00000000 ;
			15'h00003DE2 : data <= 8'b00000000 ;
			15'h00003DE3 : data <= 8'b00000000 ;
			15'h00003DE4 : data <= 8'b00000000 ;
			15'h00003DE5 : data <= 8'b00000000 ;
			15'h00003DE6 : data <= 8'b00000000 ;
			15'h00003DE7 : data <= 8'b00000000 ;
			15'h00003DE8 : data <= 8'b00000000 ;
			15'h00003DE9 : data <= 8'b00000000 ;
			15'h00003DEA : data <= 8'b00000000 ;
			15'h00003DEB : data <= 8'b00000000 ;
			15'h00003DEC : data <= 8'b00000000 ;
			15'h00003DED : data <= 8'b00000000 ;
			15'h00003DEE : data <= 8'b00000000 ;
			15'h00003DEF : data <= 8'b00000000 ;
			15'h00003DF0 : data <= 8'b00000000 ;
			15'h00003DF1 : data <= 8'b00000000 ;
			15'h00003DF2 : data <= 8'b00000000 ;
			15'h00003DF3 : data <= 8'b00000000 ;
			15'h00003DF4 : data <= 8'b00000000 ;
			15'h00003DF5 : data <= 8'b00000000 ;
			15'h00003DF6 : data <= 8'b00000000 ;
			15'h00003DF7 : data <= 8'b00000000 ;
			15'h00003DF8 : data <= 8'b00000000 ;
			15'h00003DF9 : data <= 8'b00000000 ;
			15'h00003DFA : data <= 8'b00000000 ;
			15'h00003DFB : data <= 8'b00000000 ;
			15'h00003DFC : data <= 8'b00000000 ;
			15'h00003DFD : data <= 8'b00000000 ;
			15'h00003DFE : data <= 8'b00000000 ;
			15'h00003DFF : data <= 8'b00000000 ;
			15'h00003E00 : data <= 8'b00000000 ;
			15'h00003E01 : data <= 8'b00000000 ;
			15'h00003E02 : data <= 8'b00000000 ;
			15'h00003E03 : data <= 8'b00000000 ;
			15'h00003E04 : data <= 8'b00000000 ;
			15'h00003E05 : data <= 8'b00000000 ;
			15'h00003E06 : data <= 8'b00000000 ;
			15'h00003E07 : data <= 8'b00000000 ;
			15'h00003E08 : data <= 8'b00000000 ;
			15'h00003E09 : data <= 8'b00000000 ;
			15'h00003E0A : data <= 8'b00000000 ;
			15'h00003E0B : data <= 8'b00000000 ;
			15'h00003E0C : data <= 8'b00000000 ;
			15'h00003E0D : data <= 8'b00000000 ;
			15'h00003E0E : data <= 8'b00000000 ;
			15'h00003E0F : data <= 8'b00000000 ;
			15'h00003E10 : data <= 8'b00000000 ;
			15'h00003E11 : data <= 8'b00000000 ;
			15'h00003E12 : data <= 8'b00000000 ;
			15'h00003E13 : data <= 8'b00000000 ;
			15'h00003E14 : data <= 8'b00000000 ;
			15'h00003E15 : data <= 8'b00000000 ;
			15'h00003E16 : data <= 8'b00000000 ;
			15'h00003E17 : data <= 8'b00000000 ;
			15'h00003E18 : data <= 8'b00000000 ;
			15'h00003E19 : data <= 8'b00000000 ;
			15'h00003E1A : data <= 8'b00000000 ;
			15'h00003E1B : data <= 8'b00000000 ;
			15'h00003E1C : data <= 8'b00000000 ;
			15'h00003E1D : data <= 8'b00000000 ;
			15'h00003E1E : data <= 8'b00000000 ;
			15'h00003E1F : data <= 8'b00000000 ;
			15'h00003E20 : data <= 8'b00000000 ;
			15'h00003E21 : data <= 8'b00000000 ;
			15'h00003E22 : data <= 8'b00000000 ;
			15'h00003E23 : data <= 8'b00000000 ;
			15'h00003E24 : data <= 8'b00000000 ;
			15'h00003E25 : data <= 8'b00000000 ;
			15'h00003E26 : data <= 8'b00000000 ;
			15'h00003E27 : data <= 8'b00000000 ;
			15'h00003E28 : data <= 8'b00000000 ;
			15'h00003E29 : data <= 8'b00000000 ;
			15'h00003E2A : data <= 8'b00000000 ;
			15'h00003E2B : data <= 8'b00000000 ;
			15'h00003E2C : data <= 8'b00000000 ;
			15'h00003E2D : data <= 8'b00000000 ;
			15'h00003E2E : data <= 8'b00000000 ;
			15'h00003E2F : data <= 8'b00000000 ;
			15'h00003E30 : data <= 8'b00000000 ;
			15'h00003E31 : data <= 8'b00000000 ;
			15'h00003E32 : data <= 8'b00000000 ;
			15'h00003E33 : data <= 8'b00000000 ;
			15'h00003E34 : data <= 8'b00000000 ;
			15'h00003E35 : data <= 8'b00000000 ;
			15'h00003E36 : data <= 8'b00000000 ;
			15'h00003E37 : data <= 8'b00000000 ;
			15'h00003E38 : data <= 8'b00000000 ;
			15'h00003E39 : data <= 8'b00000000 ;
			15'h00003E3A : data <= 8'b00000000 ;
			15'h00003E3B : data <= 8'b00000000 ;
			15'h00003E3C : data <= 8'b00000000 ;
			15'h00003E3D : data <= 8'b00000000 ;
			15'h00003E3E : data <= 8'b00000000 ;
			15'h00003E3F : data <= 8'b00000000 ;
			15'h00003E40 : data <= 8'b00000000 ;
			15'h00003E41 : data <= 8'b00000000 ;
			15'h00003E42 : data <= 8'b00000000 ;
			15'h00003E43 : data <= 8'b00000000 ;
			15'h00003E44 : data <= 8'b00000000 ;
			15'h00003E45 : data <= 8'b00000000 ;
			15'h00003E46 : data <= 8'b00000000 ;
			15'h00003E47 : data <= 8'b00000000 ;
			15'h00003E48 : data <= 8'b00000000 ;
			15'h00003E49 : data <= 8'b00000000 ;
			15'h00003E4A : data <= 8'b00000000 ;
			15'h00003E4B : data <= 8'b00000000 ;
			15'h00003E4C : data <= 8'b00000000 ;
			15'h00003E4D : data <= 8'b00000000 ;
			15'h00003E4E : data <= 8'b00000000 ;
			15'h00003E4F : data <= 8'b00000000 ;
			15'h00003E50 : data <= 8'b00000000 ;
			15'h00003E51 : data <= 8'b00000000 ;
			15'h00003E52 : data <= 8'b00000000 ;
			15'h00003E53 : data <= 8'b00000000 ;
			15'h00003E54 : data <= 8'b00000000 ;
			15'h00003E55 : data <= 8'b00000000 ;
			15'h00003E56 : data <= 8'b00000000 ;
			15'h00003E57 : data <= 8'b00000000 ;
			15'h00003E58 : data <= 8'b00000000 ;
			15'h00003E59 : data <= 8'b00000000 ;
			15'h00003E5A : data <= 8'b00000000 ;
			15'h00003E5B : data <= 8'b00000000 ;
			15'h00003E5C : data <= 8'b00000000 ;
			15'h00003E5D : data <= 8'b00000000 ;
			15'h00003E5E : data <= 8'b00000000 ;
			15'h00003E5F : data <= 8'b00000000 ;
			15'h00003E60 : data <= 8'b00000000 ;
			15'h00003E61 : data <= 8'b00000000 ;
			15'h00003E62 : data <= 8'b00000000 ;
			15'h00003E63 : data <= 8'b00000000 ;
			15'h00003E64 : data <= 8'b00000000 ;
			15'h00003E65 : data <= 8'b00000000 ;
			15'h00003E66 : data <= 8'b00000000 ;
			15'h00003E67 : data <= 8'b00000000 ;
			15'h00003E68 : data <= 8'b00000000 ;
			15'h00003E69 : data <= 8'b00000000 ;
			15'h00003E6A : data <= 8'b00000000 ;
			15'h00003E6B : data <= 8'b00000000 ;
			15'h00003E6C : data <= 8'b00000000 ;
			15'h00003E6D : data <= 8'b00000000 ;
			15'h00003E6E : data <= 8'b00000000 ;
			15'h00003E6F : data <= 8'b00000000 ;
			15'h00003E70 : data <= 8'b00000000 ;
			15'h00003E71 : data <= 8'b00000000 ;
			15'h00003E72 : data <= 8'b00000000 ;
			15'h00003E73 : data <= 8'b00000000 ;
			15'h00003E74 : data <= 8'b00000000 ;
			15'h00003E75 : data <= 8'b00000000 ;
			15'h00003E76 : data <= 8'b00000000 ;
			15'h00003E77 : data <= 8'b00000000 ;
			15'h00003E78 : data <= 8'b00000000 ;
			15'h00003E79 : data <= 8'b00000000 ;
			15'h00003E7A : data <= 8'b00000000 ;
			15'h00003E7B : data <= 8'b00000000 ;
			15'h00003E7C : data <= 8'b00000000 ;
			15'h00003E7D : data <= 8'b00000000 ;
			15'h00003E7E : data <= 8'b00000000 ;
			15'h00003E7F : data <= 8'b00000000 ;
			15'h00003E80 : data <= 8'b00000000 ;
			15'h00003E81 : data <= 8'b00000000 ;
			15'h00003E82 : data <= 8'b00000000 ;
			15'h00003E83 : data <= 8'b00000000 ;
			15'h00003E84 : data <= 8'b00000000 ;
			15'h00003E85 : data <= 8'b00000000 ;
			15'h00003E86 : data <= 8'b00000000 ;
			15'h00003E87 : data <= 8'b00000000 ;
			15'h00003E88 : data <= 8'b00000000 ;
			15'h00003E89 : data <= 8'b00000000 ;
			15'h00003E8A : data <= 8'b00000000 ;
			15'h00003E8B : data <= 8'b00000000 ;
			15'h00003E8C : data <= 8'b00000000 ;
			15'h00003E8D : data <= 8'b00000000 ;
			15'h00003E8E : data <= 8'b00000000 ;
			15'h00003E8F : data <= 8'b00000000 ;
			15'h00003E90 : data <= 8'b00000000 ;
			15'h00003E91 : data <= 8'b00000000 ;
			15'h00003E92 : data <= 8'b00000000 ;
			15'h00003E93 : data <= 8'b00000000 ;
			15'h00003E94 : data <= 8'b00000000 ;
			15'h00003E95 : data <= 8'b00000000 ;
			15'h00003E96 : data <= 8'b00000000 ;
			15'h00003E97 : data <= 8'b00000000 ;
			15'h00003E98 : data <= 8'b00000000 ;
			15'h00003E99 : data <= 8'b00000000 ;
			15'h00003E9A : data <= 8'b00000000 ;
			15'h00003E9B : data <= 8'b00000000 ;
			15'h00003E9C : data <= 8'b00000000 ;
			15'h00003E9D : data <= 8'b00000000 ;
			15'h00003E9E : data <= 8'b00000000 ;
			15'h00003E9F : data <= 8'b00000000 ;
			15'h00003EA0 : data <= 8'b00000000 ;
			15'h00003EA1 : data <= 8'b00000000 ;
			15'h00003EA2 : data <= 8'b00000000 ;
			15'h00003EA3 : data <= 8'b00000000 ;
			15'h00003EA4 : data <= 8'b00000000 ;
			15'h00003EA5 : data <= 8'b00000000 ;
			15'h00003EA6 : data <= 8'b00000000 ;
			15'h00003EA7 : data <= 8'b00000000 ;
			15'h00003EA8 : data <= 8'b00000000 ;
			15'h00003EA9 : data <= 8'b00000000 ;
			15'h00003EAA : data <= 8'b00000000 ;
			15'h00003EAB : data <= 8'b00000000 ;
			15'h00003EAC : data <= 8'b00000000 ;
			15'h00003EAD : data <= 8'b00000000 ;
			15'h00003EAE : data <= 8'b00000000 ;
			15'h00003EAF : data <= 8'b00000000 ;
			15'h00003EB0 : data <= 8'b00000000 ;
			15'h00003EB1 : data <= 8'b00000000 ;
			15'h00003EB2 : data <= 8'b00000000 ;
			15'h00003EB3 : data <= 8'b00000000 ;
			15'h00003EB4 : data <= 8'b00000000 ;
			15'h00003EB5 : data <= 8'b00000000 ;
			15'h00003EB6 : data <= 8'b00000000 ;
			15'h00003EB7 : data <= 8'b00000000 ;
			15'h00003EB8 : data <= 8'b00000000 ;
			15'h00003EB9 : data <= 8'b00000000 ;
			15'h00003EBA : data <= 8'b00000000 ;
			15'h00003EBB : data <= 8'b00000000 ;
			15'h00003EBC : data <= 8'b00000000 ;
			15'h00003EBD : data <= 8'b00000000 ;
			15'h00003EBE : data <= 8'b00000000 ;
			15'h00003EBF : data <= 8'b00000000 ;
			15'h00003EC0 : data <= 8'b00000000 ;
			15'h00003EC1 : data <= 8'b00000000 ;
			15'h00003EC2 : data <= 8'b00000000 ;
			15'h00003EC3 : data <= 8'b00000000 ;
			15'h00003EC4 : data <= 8'b00000000 ;
			15'h00003EC5 : data <= 8'b00000000 ;
			15'h00003EC6 : data <= 8'b00000000 ;
			15'h00003EC7 : data <= 8'b00000000 ;
			15'h00003EC8 : data <= 8'b00000000 ;
			15'h00003EC9 : data <= 8'b00000000 ;
			15'h00003ECA : data <= 8'b00000000 ;
			15'h00003ECB : data <= 8'b00000000 ;
			15'h00003ECC : data <= 8'b00000000 ;
			15'h00003ECD : data <= 8'b00000000 ;
			15'h00003ECE : data <= 8'b00000000 ;
			15'h00003ECF : data <= 8'b00000000 ;
			15'h00003ED0 : data <= 8'b00000000 ;
			15'h00003ED1 : data <= 8'b00000000 ;
			15'h00003ED2 : data <= 8'b00000000 ;
			15'h00003ED3 : data <= 8'b00000000 ;
			15'h00003ED4 : data <= 8'b00000000 ;
			15'h00003ED5 : data <= 8'b00000000 ;
			15'h00003ED6 : data <= 8'b00000000 ;
			15'h00003ED7 : data <= 8'b00000000 ;
			15'h00003ED8 : data <= 8'b00000000 ;
			15'h00003ED9 : data <= 8'b00000000 ;
			15'h00003EDA : data <= 8'b00000000 ;
			15'h00003EDB : data <= 8'b00000000 ;
			15'h00003EDC : data <= 8'b00000000 ;
			15'h00003EDD : data <= 8'b00000000 ;
			15'h00003EDE : data <= 8'b00000000 ;
			15'h00003EDF : data <= 8'b00000000 ;
			15'h00003EE0 : data <= 8'b00000000 ;
			15'h00003EE1 : data <= 8'b00000000 ;
			15'h00003EE2 : data <= 8'b00000000 ;
			15'h00003EE3 : data <= 8'b00000000 ;
			15'h00003EE4 : data <= 8'b00000000 ;
			15'h00003EE5 : data <= 8'b00000000 ;
			15'h00003EE6 : data <= 8'b00000000 ;
			15'h00003EE7 : data <= 8'b00000000 ;
			15'h00003EE8 : data <= 8'b00000000 ;
			15'h00003EE9 : data <= 8'b00000000 ;
			15'h00003EEA : data <= 8'b00000000 ;
			15'h00003EEB : data <= 8'b00000000 ;
			15'h00003EEC : data <= 8'b00000000 ;
			15'h00003EED : data <= 8'b00000000 ;
			15'h00003EEE : data <= 8'b00000000 ;
			15'h00003EEF : data <= 8'b00000000 ;
			15'h00003EF0 : data <= 8'b00000000 ;
			15'h00003EF1 : data <= 8'b00000000 ;
			15'h00003EF2 : data <= 8'b00000000 ;
			15'h00003EF3 : data <= 8'b00000000 ;
			15'h00003EF4 : data <= 8'b00000000 ;
			15'h00003EF5 : data <= 8'b00000000 ;
			15'h00003EF6 : data <= 8'b00000000 ;
			15'h00003EF7 : data <= 8'b00000000 ;
			15'h00003EF8 : data <= 8'b00000000 ;
			15'h00003EF9 : data <= 8'b00000000 ;
			15'h00003EFA : data <= 8'b00000000 ;
			15'h00003EFB : data <= 8'b00000000 ;
			15'h00003EFC : data <= 8'b00000000 ;
			15'h00003EFD : data <= 8'b00000000 ;
			15'h00003EFE : data <= 8'b00000000 ;
			15'h00003EFF : data <= 8'b00000000 ;
			15'h00003F00 : data <= 8'b00000000 ;
			15'h00003F01 : data <= 8'b00000000 ;
			15'h00003F02 : data <= 8'b00000000 ;
			15'h00003F03 : data <= 8'b00000000 ;
			15'h00003F04 : data <= 8'b00000000 ;
			15'h00003F05 : data <= 8'b00000000 ;
			15'h00003F06 : data <= 8'b00000000 ;
			15'h00003F07 : data <= 8'b00000000 ;
			15'h00003F08 : data <= 8'b00000000 ;
			15'h00003F09 : data <= 8'b00000000 ;
			15'h00003F0A : data <= 8'b00000000 ;
			15'h00003F0B : data <= 8'b00000000 ;
			15'h00003F0C : data <= 8'b00000000 ;
			15'h00003F0D : data <= 8'b00000000 ;
			15'h00003F0E : data <= 8'b00000000 ;
			15'h00003F0F : data <= 8'b00000000 ;
			15'h00003F10 : data <= 8'b00000000 ;
			15'h00003F11 : data <= 8'b00000000 ;
			15'h00003F12 : data <= 8'b00000000 ;
			15'h00003F13 : data <= 8'b00000000 ;
			15'h00003F14 : data <= 8'b00000000 ;
			15'h00003F15 : data <= 8'b00000000 ;
			15'h00003F16 : data <= 8'b00000000 ;
			15'h00003F17 : data <= 8'b00000000 ;
			15'h00003F18 : data <= 8'b00000000 ;
			15'h00003F19 : data <= 8'b00000000 ;
			15'h00003F1A : data <= 8'b00000000 ;
			15'h00003F1B : data <= 8'b00000000 ;
			15'h00003F1C : data <= 8'b00000000 ;
			15'h00003F1D : data <= 8'b00000000 ;
			15'h00003F1E : data <= 8'b00000000 ;
			15'h00003F1F : data <= 8'b00000000 ;
			15'h00003F20 : data <= 8'b00000000 ;
			15'h00003F21 : data <= 8'b00000000 ;
			15'h00003F22 : data <= 8'b00000000 ;
			15'h00003F23 : data <= 8'b00000000 ;
			15'h00003F24 : data <= 8'b00000000 ;
			15'h00003F25 : data <= 8'b00000000 ;
			15'h00003F26 : data <= 8'b00000000 ;
			15'h00003F27 : data <= 8'b00000000 ;
			15'h00003F28 : data <= 8'b00000000 ;
			15'h00003F29 : data <= 8'b00000000 ;
			15'h00003F2A : data <= 8'b00000000 ;
			15'h00003F2B : data <= 8'b00000000 ;
			15'h00003F2C : data <= 8'b00000000 ;
			15'h00003F2D : data <= 8'b00000000 ;
			15'h00003F2E : data <= 8'b00000000 ;
			15'h00003F2F : data <= 8'b00000000 ;
			15'h00003F30 : data <= 8'b00000000 ;
			15'h00003F31 : data <= 8'b00000000 ;
			15'h00003F32 : data <= 8'b00000000 ;
			15'h00003F33 : data <= 8'b00000000 ;
			15'h00003F34 : data <= 8'b00000000 ;
			15'h00003F35 : data <= 8'b00000000 ;
			15'h00003F36 : data <= 8'b00000000 ;
			15'h00003F37 : data <= 8'b00000000 ;
			15'h00003F38 : data <= 8'b00000000 ;
			15'h00003F39 : data <= 8'b00000000 ;
			15'h00003F3A : data <= 8'b00000000 ;
			15'h00003F3B : data <= 8'b00000000 ;
			15'h00003F3C : data <= 8'b00000000 ;
			15'h00003F3D : data <= 8'b00000000 ;
			15'h00003F3E : data <= 8'b00000000 ;
			15'h00003F3F : data <= 8'b00000000 ;
			15'h00003F40 : data <= 8'b00000000 ;
			15'h00003F41 : data <= 8'b00000000 ;
			15'h00003F42 : data <= 8'b00000000 ;
			15'h00003F43 : data <= 8'b00000000 ;
			15'h00003F44 : data <= 8'b00000000 ;
			15'h00003F45 : data <= 8'b00000000 ;
			15'h00003F46 : data <= 8'b00000000 ;
			15'h00003F47 : data <= 8'b00000000 ;
			15'h00003F48 : data <= 8'b00000000 ;
			15'h00003F49 : data <= 8'b00000000 ;
			15'h00003F4A : data <= 8'b00000000 ;
			15'h00003F4B : data <= 8'b00000000 ;
			15'h00003F4C : data <= 8'b00000000 ;
			15'h00003F4D : data <= 8'b00000000 ;
			15'h00003F4E : data <= 8'b00000000 ;
			15'h00003F4F : data <= 8'b00000000 ;
			15'h00003F50 : data <= 8'b00000000 ;
			15'h00003F51 : data <= 8'b00000000 ;
			15'h00003F52 : data <= 8'b00000000 ;
			15'h00003F53 : data <= 8'b00000000 ;
			15'h00003F54 : data <= 8'b00000000 ;
			15'h00003F55 : data <= 8'b00000000 ;
			15'h00003F56 : data <= 8'b00000000 ;
			15'h00003F57 : data <= 8'b00000000 ;
			15'h00003F58 : data <= 8'b00000000 ;
			15'h00003F59 : data <= 8'b00000000 ;
			15'h00003F5A : data <= 8'b00000000 ;
			15'h00003F5B : data <= 8'b00000000 ;
			15'h00003F5C : data <= 8'b00000000 ;
			15'h00003F5D : data <= 8'b00000000 ;
			15'h00003F5E : data <= 8'b00000000 ;
			15'h00003F5F : data <= 8'b00000000 ;
			15'h00003F60 : data <= 8'b00000000 ;
			15'h00003F61 : data <= 8'b00000000 ;
			15'h00003F62 : data <= 8'b00000000 ;
			15'h00003F63 : data <= 8'b00000000 ;
			15'h00003F64 : data <= 8'b00000000 ;
			15'h00003F65 : data <= 8'b00000000 ;
			15'h00003F66 : data <= 8'b00000000 ;
			15'h00003F67 : data <= 8'b00000000 ;
			15'h00003F68 : data <= 8'b00000000 ;
			15'h00003F69 : data <= 8'b00000000 ;
			15'h00003F6A : data <= 8'b00000000 ;
			15'h00003F6B : data <= 8'b00000000 ;
			15'h00003F6C : data <= 8'b00000000 ;
			15'h00003F6D : data <= 8'b00000000 ;
			15'h00003F6E : data <= 8'b00000000 ;
			15'h00003F6F : data <= 8'b00000000 ;
			15'h00003F70 : data <= 8'b00000000 ;
			15'h00003F71 : data <= 8'b00000000 ;
			15'h00003F72 : data <= 8'b00000000 ;
			15'h00003F73 : data <= 8'b00000000 ;
			15'h00003F74 : data <= 8'b00000000 ;
			15'h00003F75 : data <= 8'b00000000 ;
			15'h00003F76 : data <= 8'b00000000 ;
			15'h00003F77 : data <= 8'b00000000 ;
			15'h00003F78 : data <= 8'b00000000 ;
			15'h00003F79 : data <= 8'b00000000 ;
			15'h00003F7A : data <= 8'b00000000 ;
			15'h00003F7B : data <= 8'b00000000 ;
			15'h00003F7C : data <= 8'b00000000 ;
			15'h00003F7D : data <= 8'b00000000 ;
			15'h00003F7E : data <= 8'b00000000 ;
			15'h00003F7F : data <= 8'b00000000 ;
			15'h00003F80 : data <= 8'b00000000 ;
			15'h00003F81 : data <= 8'b00000000 ;
			15'h00003F82 : data <= 8'b00000000 ;
			15'h00003F83 : data <= 8'b00000000 ;
			15'h00003F84 : data <= 8'b00000000 ;
			15'h00003F85 : data <= 8'b00000000 ;
			15'h00003F86 : data <= 8'b00000000 ;
			15'h00003F87 : data <= 8'b00000000 ;
			15'h00003F88 : data <= 8'b00000000 ;
			15'h00003F89 : data <= 8'b00000000 ;
			15'h00003F8A : data <= 8'b00000000 ;
			15'h00003F8B : data <= 8'b00000000 ;
			15'h00003F8C : data <= 8'b00000000 ;
			15'h00003F8D : data <= 8'b00000000 ;
			15'h00003F8E : data <= 8'b00000000 ;
			15'h00003F8F : data <= 8'b00000000 ;
			15'h00003F90 : data <= 8'b00000000 ;
			15'h00003F91 : data <= 8'b00000000 ;
			15'h00003F92 : data <= 8'b00000000 ;
			15'h00003F93 : data <= 8'b00000000 ;
			15'h00003F94 : data <= 8'b00000000 ;
			15'h00003F95 : data <= 8'b00000000 ;
			15'h00003F96 : data <= 8'b00000000 ;
			15'h00003F97 : data <= 8'b00000000 ;
			15'h00003F98 : data <= 8'b00000000 ;
			15'h00003F99 : data <= 8'b00000000 ;
			15'h00003F9A : data <= 8'b00000000 ;
			15'h00003F9B : data <= 8'b00000000 ;
			15'h00003F9C : data <= 8'b00000000 ;
			15'h00003F9D : data <= 8'b00000000 ;
			15'h00003F9E : data <= 8'b00000000 ;
			15'h00003F9F : data <= 8'b00000000 ;
			15'h00003FA0 : data <= 8'b00000000 ;
			15'h00003FA1 : data <= 8'b00000000 ;
			15'h00003FA2 : data <= 8'b00000000 ;
			15'h00003FA3 : data <= 8'b00000000 ;
			15'h00003FA4 : data <= 8'b00000000 ;
			15'h00003FA5 : data <= 8'b00000000 ;
			15'h00003FA6 : data <= 8'b00000000 ;
			15'h00003FA7 : data <= 8'b00000000 ;
			15'h00003FA8 : data <= 8'b00000000 ;
			15'h00003FA9 : data <= 8'b00000000 ;
			15'h00003FAA : data <= 8'b00000000 ;
			15'h00003FAB : data <= 8'b00000000 ;
			15'h00003FAC : data <= 8'b00000000 ;
			15'h00003FAD : data <= 8'b00000000 ;
			15'h00003FAE : data <= 8'b00000000 ;
			15'h00003FAF : data <= 8'b00000000 ;
			15'h00003FB0 : data <= 8'b00000000 ;
			15'h00003FB1 : data <= 8'b00000000 ;
			15'h00003FB2 : data <= 8'b00000000 ;
			15'h00003FB3 : data <= 8'b00000000 ;
			15'h00003FB4 : data <= 8'b00000000 ;
			15'h00003FB5 : data <= 8'b00000000 ;
			15'h00003FB6 : data <= 8'b00000000 ;
			15'h00003FB7 : data <= 8'b00000000 ;
			15'h00003FB8 : data <= 8'b00000000 ;
			15'h00003FB9 : data <= 8'b00000000 ;
			15'h00003FBA : data <= 8'b00000000 ;
			15'h00003FBB : data <= 8'b00000000 ;
			15'h00003FBC : data <= 8'b00000000 ;
			15'h00003FBD : data <= 8'b00000000 ;
			15'h00003FBE : data <= 8'b00000000 ;
			15'h00003FBF : data <= 8'b00000000 ;
			15'h00003FC0 : data <= 8'b00000000 ;
			15'h00003FC1 : data <= 8'b00000000 ;
			15'h00003FC2 : data <= 8'b00000000 ;
			15'h00003FC3 : data <= 8'b00000000 ;
			15'h00003FC4 : data <= 8'b00000000 ;
			15'h00003FC5 : data <= 8'b00000000 ;
			15'h00003FC6 : data <= 8'b00000000 ;
			15'h00003FC7 : data <= 8'b00000000 ;
			15'h00003FC8 : data <= 8'b00000000 ;
			15'h00003FC9 : data <= 8'b00000000 ;
			15'h00003FCA : data <= 8'b00000000 ;
			15'h00003FCB : data <= 8'b00000000 ;
			15'h00003FCC : data <= 8'b00000000 ;
			15'h00003FCD : data <= 8'b00000000 ;
			15'h00003FCE : data <= 8'b00000000 ;
			15'h00003FCF : data <= 8'b00000000 ;
			15'h00003FD0 : data <= 8'b00000000 ;
			15'h00003FD1 : data <= 8'b00000000 ;
			15'h00003FD2 : data <= 8'b00000000 ;
			15'h00003FD3 : data <= 8'b00000000 ;
			15'h00003FD4 : data <= 8'b00000000 ;
			15'h00003FD5 : data <= 8'b00000000 ;
			15'h00003FD6 : data <= 8'b00000000 ;
			15'h00003FD7 : data <= 8'b00000000 ;
			15'h00003FD8 : data <= 8'b00000000 ;
			15'h00003FD9 : data <= 8'b00000000 ;
			15'h00003FDA : data <= 8'b00000000 ;
			15'h00003FDB : data <= 8'b00000000 ;
			15'h00003FDC : data <= 8'b00000000 ;
			15'h00003FDD : data <= 8'b00000000 ;
			15'h00003FDE : data <= 8'b00000000 ;
			15'h00003FDF : data <= 8'b00000000 ;
			15'h00003FE0 : data <= 8'b00000000 ;
			15'h00003FE1 : data <= 8'b00000000 ;
			15'h00003FE2 : data <= 8'b00000000 ;
			15'h00003FE3 : data <= 8'b00000000 ;
			15'h00003FE4 : data <= 8'b00000000 ;
			15'h00003FE5 : data <= 8'b00000000 ;
			15'h00003FE6 : data <= 8'b00000000 ;
			15'h00003FE7 : data <= 8'b00000000 ;
			15'h00003FE8 : data <= 8'b00000000 ;
			15'h00003FE9 : data <= 8'b00000000 ;
			15'h00003FEA : data <= 8'b00000000 ;
			15'h00003FEB : data <= 8'b00000000 ;
			15'h00003FEC : data <= 8'b00000000 ;
			15'h00003FED : data <= 8'b00000000 ;
			15'h00003FEE : data <= 8'b00000000 ;
			15'h00003FEF : data <= 8'b00000000 ;
			15'h00003FF0 : data <= 8'b00000000 ;
			15'h00003FF1 : data <= 8'b00000000 ;
			15'h00003FF2 : data <= 8'b00000000 ;
			15'h00003FF3 : data <= 8'b00000000 ;
			15'h00003FF4 : data <= 8'b00000000 ;
			15'h00003FF5 : data <= 8'b00000000 ;
			15'h00003FF6 : data <= 8'b00000000 ;
			15'h00003FF7 : data <= 8'b00000000 ;
			15'h00003FF8 : data <= 8'b00000000 ;
			15'h00003FF9 : data <= 8'b00000000 ;
			15'h00003FFA : data <= 8'b00000000 ;
			15'h00003FFB : data <= 8'b00000000 ;
			15'h00003FFC : data <= 8'b00000000 ;
			15'h00003FFD : data <= 8'b00000000 ;
			15'h00003FFE : data <= 8'b00000000 ;
			15'h00003FFF : data <= 8'b00000000 ;
			15'h00004000 : data <= 8'b00000000 ;
			15'h00004001 : data <= 8'b00000000 ;
			15'h00004002 : data <= 8'b00000000 ;
			15'h00004003 : data <= 8'b00000000 ;
			15'h00004004 : data <= 8'b00000000 ;
			15'h00004005 : data <= 8'b00000000 ;
			15'h00004006 : data <= 8'b00000000 ;
			15'h00004007 : data <= 8'b00000000 ;
			15'h00004008 : data <= 8'b00000000 ;
			15'h00004009 : data <= 8'b00000000 ;
			15'h0000400A : data <= 8'b00000000 ;
			15'h0000400B : data <= 8'b00000000 ;
			15'h0000400C : data <= 8'b00000000 ;
			15'h0000400D : data <= 8'b00000000 ;
			15'h0000400E : data <= 8'b00000000 ;
			15'h0000400F : data <= 8'b00000000 ;
			15'h00004010 : data <= 8'b00000000 ;
			15'h00004011 : data <= 8'b00000000 ;
			15'h00004012 : data <= 8'b00000000 ;
			15'h00004013 : data <= 8'b00000000 ;
			15'h00004014 : data <= 8'b00000000 ;
			15'h00004015 : data <= 8'b00000000 ;
			15'h00004016 : data <= 8'b00000000 ;
			15'h00004017 : data <= 8'b00000000 ;
			15'h00004018 : data <= 8'b00000000 ;
			15'h00004019 : data <= 8'b00000000 ;
			15'h0000401A : data <= 8'b00000000 ;
			15'h0000401B : data <= 8'b00000000 ;
			15'h0000401C : data <= 8'b00000000 ;
			15'h0000401D : data <= 8'b00000000 ;
			15'h0000401E : data <= 8'b00000000 ;
			15'h0000401F : data <= 8'b00000000 ;
			15'h00004020 : data <= 8'b00000000 ;
			15'h00004021 : data <= 8'b00000000 ;
			15'h00004022 : data <= 8'b00000000 ;
			15'h00004023 : data <= 8'b00000000 ;
			15'h00004024 : data <= 8'b00000000 ;
			15'h00004025 : data <= 8'b00000000 ;
			15'h00004026 : data <= 8'b00000000 ;
			15'h00004027 : data <= 8'b00000000 ;
			15'h00004028 : data <= 8'b00000000 ;
			15'h00004029 : data <= 8'b00000000 ;
			15'h0000402A : data <= 8'b00000000 ;
			15'h0000402B : data <= 8'b00000000 ;
			15'h0000402C : data <= 8'b00000000 ;
			15'h0000402D : data <= 8'b00000000 ;
			15'h0000402E : data <= 8'b00000000 ;
			15'h0000402F : data <= 8'b00000000 ;
			15'h00004030 : data <= 8'b00000000 ;
			15'h00004031 : data <= 8'b00000000 ;
			15'h00004032 : data <= 8'b00000000 ;
			15'h00004033 : data <= 8'b00000000 ;
			15'h00004034 : data <= 8'b00000000 ;
			15'h00004035 : data <= 8'b00000000 ;
			15'h00004036 : data <= 8'b00000000 ;
			15'h00004037 : data <= 8'b00000000 ;
			15'h00004038 : data <= 8'b00000000 ;
			15'h00004039 : data <= 8'b00000000 ;
			15'h0000403A : data <= 8'b00000000 ;
			15'h0000403B : data <= 8'b00000000 ;
			15'h0000403C : data <= 8'b00000000 ;
			15'h0000403D : data <= 8'b00000000 ;
			15'h0000403E : data <= 8'b00000000 ;
			15'h0000403F : data <= 8'b00000000 ;
			15'h00004040 : data <= 8'b00000000 ;
			15'h00004041 : data <= 8'b00000000 ;
			15'h00004042 : data <= 8'b00000000 ;
			15'h00004043 : data <= 8'b00000000 ;
			15'h00004044 : data <= 8'b00000000 ;
			15'h00004045 : data <= 8'b00000000 ;
			15'h00004046 : data <= 8'b00000000 ;
			15'h00004047 : data <= 8'b00000000 ;
			15'h00004048 : data <= 8'b00000000 ;
			15'h00004049 : data <= 8'b00000000 ;
			15'h0000404A : data <= 8'b00000000 ;
			15'h0000404B : data <= 8'b00000000 ;
			15'h0000404C : data <= 8'b00000000 ;
			15'h0000404D : data <= 8'b00000000 ;
			15'h0000404E : data <= 8'b00000000 ;
			15'h0000404F : data <= 8'b00000000 ;
			15'h00004050 : data <= 8'b00000000 ;
			15'h00004051 : data <= 8'b00000000 ;
			15'h00004052 : data <= 8'b00000000 ;
			15'h00004053 : data <= 8'b00000000 ;
			15'h00004054 : data <= 8'b00000000 ;
			15'h00004055 : data <= 8'b00000000 ;
			15'h00004056 : data <= 8'b00000000 ;
			15'h00004057 : data <= 8'b00000000 ;
			15'h00004058 : data <= 8'b00000000 ;
			15'h00004059 : data <= 8'b00000000 ;
			15'h0000405A : data <= 8'b00000000 ;
			15'h0000405B : data <= 8'b00000000 ;
			15'h0000405C : data <= 8'b00000000 ;
			15'h0000405D : data <= 8'b00000000 ;
			15'h0000405E : data <= 8'b00000000 ;
			15'h0000405F : data <= 8'b00000000 ;
			15'h00004060 : data <= 8'b00000000 ;
			15'h00004061 : data <= 8'b00000000 ;
			15'h00004062 : data <= 8'b00000000 ;
			15'h00004063 : data <= 8'b00000000 ;
			15'h00004064 : data <= 8'b00000000 ;
			15'h00004065 : data <= 8'b00000000 ;
			15'h00004066 : data <= 8'b00000000 ;
			15'h00004067 : data <= 8'b00000000 ;
			15'h00004068 : data <= 8'b00000000 ;
			15'h00004069 : data <= 8'b00000000 ;
			15'h0000406A : data <= 8'b00000000 ;
			15'h0000406B : data <= 8'b00000000 ;
			15'h0000406C : data <= 8'b00000000 ;
			15'h0000406D : data <= 8'b00000000 ;
			15'h0000406E : data <= 8'b00000000 ;
			15'h0000406F : data <= 8'b00000000 ;
			15'h00004070 : data <= 8'b00000000 ;
			15'h00004071 : data <= 8'b00000000 ;
			15'h00004072 : data <= 8'b00000000 ;
			15'h00004073 : data <= 8'b00000000 ;
			15'h00004074 : data <= 8'b00000000 ;
			15'h00004075 : data <= 8'b00000000 ;
			15'h00004076 : data <= 8'b00000000 ;
			15'h00004077 : data <= 8'b00000000 ;
			15'h00004078 : data <= 8'b00000000 ;
			15'h00004079 : data <= 8'b00000000 ;
			15'h0000407A : data <= 8'b00000000 ;
			15'h0000407B : data <= 8'b00000000 ;
			15'h0000407C : data <= 8'b00000000 ;
			15'h0000407D : data <= 8'b00000000 ;
			15'h0000407E : data <= 8'b00000000 ;
			15'h0000407F : data <= 8'b00000000 ;
			15'h00004080 : data <= 8'b00000000 ;
			15'h00004081 : data <= 8'b00000000 ;
			15'h00004082 : data <= 8'b00000000 ;
			15'h00004083 : data <= 8'b00000000 ;
			15'h00004084 : data <= 8'b00000000 ;
			15'h00004085 : data <= 8'b00000000 ;
			15'h00004086 : data <= 8'b00000000 ;
			15'h00004087 : data <= 8'b00000000 ;
			15'h00004088 : data <= 8'b00000000 ;
			15'h00004089 : data <= 8'b00000000 ;
			15'h0000408A : data <= 8'b00000000 ;
			15'h0000408B : data <= 8'b00000000 ;
			15'h0000408C : data <= 8'b00000000 ;
			15'h0000408D : data <= 8'b00000000 ;
			15'h0000408E : data <= 8'b00000000 ;
			15'h0000408F : data <= 8'b00000000 ;
			15'h00004090 : data <= 8'b00000000 ;
			15'h00004091 : data <= 8'b00000000 ;
			15'h00004092 : data <= 8'b00000000 ;
			15'h00004093 : data <= 8'b00000000 ;
			15'h00004094 : data <= 8'b00000000 ;
			15'h00004095 : data <= 8'b00000000 ;
			15'h00004096 : data <= 8'b00000000 ;
			15'h00004097 : data <= 8'b00000000 ;
			15'h00004098 : data <= 8'b00000000 ;
			15'h00004099 : data <= 8'b00000000 ;
			15'h0000409A : data <= 8'b00000000 ;
			15'h0000409B : data <= 8'b00000000 ;
			15'h0000409C : data <= 8'b00000000 ;
			15'h0000409D : data <= 8'b00000000 ;
			15'h0000409E : data <= 8'b00000000 ;
			15'h0000409F : data <= 8'b00000000 ;
			15'h000040A0 : data <= 8'b00000000 ;
			15'h000040A1 : data <= 8'b00000000 ;
			15'h000040A2 : data <= 8'b00000000 ;
			15'h000040A3 : data <= 8'b00000000 ;
			15'h000040A4 : data <= 8'b00000000 ;
			15'h000040A5 : data <= 8'b00000000 ;
			15'h000040A6 : data <= 8'b00000000 ;
			15'h000040A7 : data <= 8'b00000000 ;
			15'h000040A8 : data <= 8'b00000000 ;
			15'h000040A9 : data <= 8'b00000000 ;
			15'h000040AA : data <= 8'b00000000 ;
			15'h000040AB : data <= 8'b00000000 ;
			15'h000040AC : data <= 8'b00000000 ;
			15'h000040AD : data <= 8'b00000000 ;
			15'h000040AE : data <= 8'b00000000 ;
			15'h000040AF : data <= 8'b00000000 ;
			15'h000040B0 : data <= 8'b00000000 ;
			15'h000040B1 : data <= 8'b00000000 ;
			15'h000040B2 : data <= 8'b00000000 ;
			15'h000040B3 : data <= 8'b00000000 ;
			15'h000040B4 : data <= 8'b00000000 ;
			15'h000040B5 : data <= 8'b00000000 ;
			15'h000040B6 : data <= 8'b00000000 ;
			15'h000040B7 : data <= 8'b00000000 ;
			15'h000040B8 : data <= 8'b00000000 ;
			15'h000040B9 : data <= 8'b00000000 ;
			15'h000040BA : data <= 8'b00000000 ;
			15'h000040BB : data <= 8'b00000000 ;
			15'h000040BC : data <= 8'b00000000 ;
			15'h000040BD : data <= 8'b00000000 ;
			15'h000040BE : data <= 8'b00000000 ;
			15'h000040BF : data <= 8'b00000000 ;
			15'h000040C0 : data <= 8'b00000000 ;
			15'h000040C1 : data <= 8'b00000000 ;
			15'h000040C2 : data <= 8'b00000000 ;
			15'h000040C3 : data <= 8'b00000000 ;
			15'h000040C4 : data <= 8'b00000000 ;
			15'h000040C5 : data <= 8'b00000000 ;
			15'h000040C6 : data <= 8'b00000000 ;
			15'h000040C7 : data <= 8'b00000000 ;
			15'h000040C8 : data <= 8'b00000000 ;
			15'h000040C9 : data <= 8'b00000000 ;
			15'h000040CA : data <= 8'b00000000 ;
			15'h000040CB : data <= 8'b00000000 ;
			15'h000040CC : data <= 8'b00000000 ;
			15'h000040CD : data <= 8'b00000000 ;
			15'h000040CE : data <= 8'b00000000 ;
			15'h000040CF : data <= 8'b00000000 ;
			15'h000040D0 : data <= 8'b00000000 ;
			15'h000040D1 : data <= 8'b00000000 ;
			15'h000040D2 : data <= 8'b00000000 ;
			15'h000040D3 : data <= 8'b00000000 ;
			15'h000040D4 : data <= 8'b00000000 ;
			15'h000040D5 : data <= 8'b00000000 ;
			15'h000040D6 : data <= 8'b00000000 ;
			15'h000040D7 : data <= 8'b00000000 ;
			15'h000040D8 : data <= 8'b00000000 ;
			15'h000040D9 : data <= 8'b00000000 ;
			15'h000040DA : data <= 8'b00000000 ;
			15'h000040DB : data <= 8'b00000000 ;
			15'h000040DC : data <= 8'b00000000 ;
			15'h000040DD : data <= 8'b00000000 ;
			15'h000040DE : data <= 8'b00000000 ;
			15'h000040DF : data <= 8'b00000000 ;
			15'h000040E0 : data <= 8'b00000000 ;
			15'h000040E1 : data <= 8'b00000000 ;
			15'h000040E2 : data <= 8'b00000000 ;
			15'h000040E3 : data <= 8'b00000000 ;
			15'h000040E4 : data <= 8'b00000000 ;
			15'h000040E5 : data <= 8'b00000000 ;
			15'h000040E6 : data <= 8'b00000000 ;
			15'h000040E7 : data <= 8'b00000000 ;
			15'h000040E8 : data <= 8'b00000000 ;
			15'h000040E9 : data <= 8'b00000000 ;
			15'h000040EA : data <= 8'b00000000 ;
			15'h000040EB : data <= 8'b00000000 ;
			15'h000040EC : data <= 8'b00000000 ;
			15'h000040ED : data <= 8'b00000000 ;
			15'h000040EE : data <= 8'b00000000 ;
			15'h000040EF : data <= 8'b00000000 ;
			15'h000040F0 : data <= 8'b00000000 ;
			15'h000040F1 : data <= 8'b00000000 ;
			15'h000040F2 : data <= 8'b00000000 ;
			15'h000040F3 : data <= 8'b00000000 ;
			15'h000040F4 : data <= 8'b00000000 ;
			15'h000040F5 : data <= 8'b00000000 ;
			15'h000040F6 : data <= 8'b00000000 ;
			15'h000040F7 : data <= 8'b00000000 ;
			15'h000040F8 : data <= 8'b00000000 ;
			15'h000040F9 : data <= 8'b00000000 ;
			15'h000040FA : data <= 8'b00000000 ;
			15'h000040FB : data <= 8'b00000000 ;
			15'h000040FC : data <= 8'b00000000 ;
			15'h000040FD : data <= 8'b00000000 ;
			15'h000040FE : data <= 8'b00000000 ;
			15'h000040FF : data <= 8'b00000000 ;
			15'h00004100 : data <= 8'b00000000 ;
			15'h00004101 : data <= 8'b00000000 ;
			15'h00004102 : data <= 8'b00000000 ;
			15'h00004103 : data <= 8'b00000000 ;
			15'h00004104 : data <= 8'b00000000 ;
			15'h00004105 : data <= 8'b00000000 ;
			15'h00004106 : data <= 8'b00000000 ;
			15'h00004107 : data <= 8'b00000000 ;
			15'h00004108 : data <= 8'b00000000 ;
			15'h00004109 : data <= 8'b00000000 ;
			15'h0000410A : data <= 8'b00000000 ;
			15'h0000410B : data <= 8'b00000000 ;
			15'h0000410C : data <= 8'b00000000 ;
			15'h0000410D : data <= 8'b00000000 ;
			15'h0000410E : data <= 8'b00000000 ;
			15'h0000410F : data <= 8'b00000000 ;
			15'h00004110 : data <= 8'b00000000 ;
			15'h00004111 : data <= 8'b00000000 ;
			15'h00004112 : data <= 8'b00000000 ;
			15'h00004113 : data <= 8'b00000000 ;
			15'h00004114 : data <= 8'b00000000 ;
			15'h00004115 : data <= 8'b00000000 ;
			15'h00004116 : data <= 8'b00000000 ;
			15'h00004117 : data <= 8'b00000000 ;
			15'h00004118 : data <= 8'b00000000 ;
			15'h00004119 : data <= 8'b00000000 ;
			15'h0000411A : data <= 8'b00000000 ;
			15'h0000411B : data <= 8'b00000000 ;
			15'h0000411C : data <= 8'b00000000 ;
			15'h0000411D : data <= 8'b00000000 ;
			15'h0000411E : data <= 8'b00000000 ;
			15'h0000411F : data <= 8'b00000000 ;
			15'h00004120 : data <= 8'b00000000 ;
			15'h00004121 : data <= 8'b00000000 ;
			15'h00004122 : data <= 8'b00000000 ;
			15'h00004123 : data <= 8'b00000000 ;
			15'h00004124 : data <= 8'b00000000 ;
			15'h00004125 : data <= 8'b00000000 ;
			15'h00004126 : data <= 8'b00000000 ;
			15'h00004127 : data <= 8'b00000000 ;
			15'h00004128 : data <= 8'b00000000 ;
			15'h00004129 : data <= 8'b00000000 ;
			15'h0000412A : data <= 8'b00000000 ;
			15'h0000412B : data <= 8'b00000000 ;
			15'h0000412C : data <= 8'b00000000 ;
			15'h0000412D : data <= 8'b00000000 ;
			15'h0000412E : data <= 8'b00000000 ;
			15'h0000412F : data <= 8'b00000000 ;
			15'h00004130 : data <= 8'b00000000 ;
			15'h00004131 : data <= 8'b00000000 ;
			15'h00004132 : data <= 8'b00000000 ;
			15'h00004133 : data <= 8'b00000000 ;
			15'h00004134 : data <= 8'b00000000 ;
			15'h00004135 : data <= 8'b00000000 ;
			15'h00004136 : data <= 8'b00000000 ;
			15'h00004137 : data <= 8'b00000000 ;
			15'h00004138 : data <= 8'b00000000 ;
			15'h00004139 : data <= 8'b00000000 ;
			15'h0000413A : data <= 8'b00000000 ;
			15'h0000413B : data <= 8'b00000000 ;
			15'h0000413C : data <= 8'b00000000 ;
			15'h0000413D : data <= 8'b00000000 ;
			15'h0000413E : data <= 8'b00000000 ;
			15'h0000413F : data <= 8'b00000000 ;
			15'h00004140 : data <= 8'b00000000 ;
			15'h00004141 : data <= 8'b00000000 ;
			15'h00004142 : data <= 8'b00000000 ;
			15'h00004143 : data <= 8'b00000000 ;
			15'h00004144 : data <= 8'b00000000 ;
			15'h00004145 : data <= 8'b00000000 ;
			15'h00004146 : data <= 8'b00000000 ;
			15'h00004147 : data <= 8'b00000000 ;
			15'h00004148 : data <= 8'b00000000 ;
			15'h00004149 : data <= 8'b00000000 ;
			15'h0000414A : data <= 8'b00000000 ;
			15'h0000414B : data <= 8'b00000000 ;
			15'h0000414C : data <= 8'b00000000 ;
			15'h0000414D : data <= 8'b00000000 ;
			15'h0000414E : data <= 8'b00000000 ;
			15'h0000414F : data <= 8'b00000000 ;
			15'h00004150 : data <= 8'b00000000 ;
			15'h00004151 : data <= 8'b00000000 ;
			15'h00004152 : data <= 8'b00000000 ;
			15'h00004153 : data <= 8'b00000000 ;
			15'h00004154 : data <= 8'b00000000 ;
			15'h00004155 : data <= 8'b00000000 ;
			15'h00004156 : data <= 8'b00000000 ;
			15'h00004157 : data <= 8'b00000000 ;
			15'h00004158 : data <= 8'b00000000 ;
			15'h00004159 : data <= 8'b00000000 ;
			15'h0000415A : data <= 8'b00000000 ;
			15'h0000415B : data <= 8'b00000000 ;
			15'h0000415C : data <= 8'b00000000 ;
			15'h0000415D : data <= 8'b00000000 ;
			15'h0000415E : data <= 8'b00000000 ;
			15'h0000415F : data <= 8'b00000000 ;
			15'h00004160 : data <= 8'b00000000 ;
			15'h00004161 : data <= 8'b00000000 ;
			15'h00004162 : data <= 8'b00000000 ;
			15'h00004163 : data <= 8'b00000000 ;
			15'h00004164 : data <= 8'b00000000 ;
			15'h00004165 : data <= 8'b00000000 ;
			15'h00004166 : data <= 8'b00000000 ;
			15'h00004167 : data <= 8'b00000000 ;
			15'h00004168 : data <= 8'b00000000 ;
			15'h00004169 : data <= 8'b00000000 ;
			15'h0000416A : data <= 8'b00000000 ;
			15'h0000416B : data <= 8'b00000000 ;
			15'h0000416C : data <= 8'b00000000 ;
			15'h0000416D : data <= 8'b00000000 ;
			15'h0000416E : data <= 8'b00000000 ;
			15'h0000416F : data <= 8'b00000000 ;
			15'h00004170 : data <= 8'b00000000 ;
			15'h00004171 : data <= 8'b00000000 ;
			15'h00004172 : data <= 8'b00000000 ;
			15'h00004173 : data <= 8'b00000000 ;
			15'h00004174 : data <= 8'b00000000 ;
			15'h00004175 : data <= 8'b00000000 ;
			15'h00004176 : data <= 8'b00000000 ;
			15'h00004177 : data <= 8'b00000000 ;
			15'h00004178 : data <= 8'b00000000 ;
			15'h00004179 : data <= 8'b00000000 ;
			15'h0000417A : data <= 8'b00000000 ;
			15'h0000417B : data <= 8'b00000000 ;
			15'h0000417C : data <= 8'b00000000 ;
			15'h0000417D : data <= 8'b00000000 ;
			15'h0000417E : data <= 8'b00000000 ;
			15'h0000417F : data <= 8'b00000000 ;
			15'h00004180 : data <= 8'b00000000 ;
			15'h00004181 : data <= 8'b00000000 ;
			15'h00004182 : data <= 8'b00000000 ;
			15'h00004183 : data <= 8'b00000000 ;
			15'h00004184 : data <= 8'b00000000 ;
			15'h00004185 : data <= 8'b00000000 ;
			15'h00004186 : data <= 8'b00000000 ;
			15'h00004187 : data <= 8'b00000000 ;
			15'h00004188 : data <= 8'b00000000 ;
			15'h00004189 : data <= 8'b00000000 ;
			15'h0000418A : data <= 8'b00000000 ;
			15'h0000418B : data <= 8'b00000000 ;
			15'h0000418C : data <= 8'b00000000 ;
			15'h0000418D : data <= 8'b00000000 ;
			15'h0000418E : data <= 8'b00000000 ;
			15'h0000418F : data <= 8'b00000000 ;
			15'h00004190 : data <= 8'b00000000 ;
			15'h00004191 : data <= 8'b00000000 ;
			15'h00004192 : data <= 8'b00000000 ;
			15'h00004193 : data <= 8'b00000000 ;
			15'h00004194 : data <= 8'b00000000 ;
			15'h00004195 : data <= 8'b00000000 ;
			15'h00004196 : data <= 8'b00000000 ;
			15'h00004197 : data <= 8'b00000000 ;
			15'h00004198 : data <= 8'b00000000 ;
			15'h00004199 : data <= 8'b00000000 ;
			15'h0000419A : data <= 8'b00000000 ;
			15'h0000419B : data <= 8'b00000000 ;
			15'h0000419C : data <= 8'b00000000 ;
			15'h0000419D : data <= 8'b00000000 ;
			15'h0000419E : data <= 8'b00000000 ;
			15'h0000419F : data <= 8'b00000000 ;
			15'h000041A0 : data <= 8'b00000000 ;
			15'h000041A1 : data <= 8'b00000000 ;
			15'h000041A2 : data <= 8'b00000000 ;
			15'h000041A3 : data <= 8'b00000000 ;
			15'h000041A4 : data <= 8'b00000000 ;
			15'h000041A5 : data <= 8'b00000000 ;
			15'h000041A6 : data <= 8'b00000000 ;
			15'h000041A7 : data <= 8'b00000000 ;
			15'h000041A8 : data <= 8'b00000000 ;
			15'h000041A9 : data <= 8'b00000000 ;
			15'h000041AA : data <= 8'b00000000 ;
			15'h000041AB : data <= 8'b00000000 ;
			15'h000041AC : data <= 8'b00000000 ;
			15'h000041AD : data <= 8'b00000000 ;
			15'h000041AE : data <= 8'b00000000 ;
			15'h000041AF : data <= 8'b00000000 ;
			15'h000041B0 : data <= 8'b00000000 ;
			15'h000041B1 : data <= 8'b00000000 ;
			15'h000041B2 : data <= 8'b00000000 ;
			15'h000041B3 : data <= 8'b00000000 ;
			15'h000041B4 : data <= 8'b00000000 ;
			15'h000041B5 : data <= 8'b00000000 ;
			15'h000041B6 : data <= 8'b00000000 ;
			15'h000041B7 : data <= 8'b00000000 ;
			15'h000041B8 : data <= 8'b00000000 ;
			15'h000041B9 : data <= 8'b00000000 ;
			15'h000041BA : data <= 8'b00000000 ;
			15'h000041BB : data <= 8'b00000000 ;
			15'h000041BC : data <= 8'b00000000 ;
			15'h000041BD : data <= 8'b00000000 ;
			15'h000041BE : data <= 8'b00000000 ;
			15'h000041BF : data <= 8'b00000000 ;
			15'h000041C0 : data <= 8'b00000000 ;
			15'h000041C1 : data <= 8'b00000000 ;
			15'h000041C2 : data <= 8'b00000000 ;
			15'h000041C3 : data <= 8'b00000000 ;
			15'h000041C4 : data <= 8'b00000000 ;
			15'h000041C5 : data <= 8'b00000000 ;
			15'h000041C6 : data <= 8'b00000000 ;
			15'h000041C7 : data <= 8'b00000000 ;
			15'h000041C8 : data <= 8'b00000000 ;
			15'h000041C9 : data <= 8'b00000000 ;
			15'h000041CA : data <= 8'b00000000 ;
			15'h000041CB : data <= 8'b00000000 ;
			15'h000041CC : data <= 8'b00000000 ;
			15'h000041CD : data <= 8'b00000000 ;
			15'h000041CE : data <= 8'b00000000 ;
			15'h000041CF : data <= 8'b00000000 ;
			15'h000041D0 : data <= 8'b00000000 ;
			15'h000041D1 : data <= 8'b00000000 ;
			15'h000041D2 : data <= 8'b00000000 ;
			15'h000041D3 : data <= 8'b00000000 ;
			15'h000041D4 : data <= 8'b00000000 ;
			15'h000041D5 : data <= 8'b00000000 ;
			15'h000041D6 : data <= 8'b00000000 ;
			15'h000041D7 : data <= 8'b00000000 ;
			15'h000041D8 : data <= 8'b00000000 ;
			15'h000041D9 : data <= 8'b00000000 ;
			15'h000041DA : data <= 8'b00000000 ;
			15'h000041DB : data <= 8'b00000000 ;
			15'h000041DC : data <= 8'b00000000 ;
			15'h000041DD : data <= 8'b00000000 ;
			15'h000041DE : data <= 8'b00000000 ;
			15'h000041DF : data <= 8'b00000000 ;
			15'h000041E0 : data <= 8'b00000000 ;
			15'h000041E1 : data <= 8'b00000000 ;
			15'h000041E2 : data <= 8'b00000000 ;
			15'h000041E3 : data <= 8'b00000000 ;
			15'h000041E4 : data <= 8'b00000000 ;
			15'h000041E5 : data <= 8'b00000000 ;
			15'h000041E6 : data <= 8'b00000000 ;
			15'h000041E7 : data <= 8'b00000000 ;
			15'h000041E8 : data <= 8'b00000000 ;
			15'h000041E9 : data <= 8'b00000000 ;
			15'h000041EA : data <= 8'b00000000 ;
			15'h000041EB : data <= 8'b00000000 ;
			15'h000041EC : data <= 8'b00000000 ;
			15'h000041ED : data <= 8'b00000000 ;
			15'h000041EE : data <= 8'b00000000 ;
			15'h000041EF : data <= 8'b00000000 ;
			15'h000041F0 : data <= 8'b00000000 ;
			15'h000041F1 : data <= 8'b00000000 ;
			15'h000041F2 : data <= 8'b00000000 ;
			15'h000041F3 : data <= 8'b00000000 ;
			15'h000041F4 : data <= 8'b00000000 ;
			15'h000041F5 : data <= 8'b00000000 ;
			15'h000041F6 : data <= 8'b00000000 ;
			15'h000041F7 : data <= 8'b00000000 ;
			15'h000041F8 : data <= 8'b00000000 ;
			15'h000041F9 : data <= 8'b00000000 ;
			15'h000041FA : data <= 8'b00000000 ;
			15'h000041FB : data <= 8'b00000000 ;
			15'h000041FC : data <= 8'b00000000 ;
			15'h000041FD : data <= 8'b00000000 ;
			15'h000041FE : data <= 8'b00000000 ;
			15'h000041FF : data <= 8'b00000000 ;
			15'h00004200 : data <= 8'b00000000 ;
			15'h00004201 : data <= 8'b00000000 ;
			15'h00004202 : data <= 8'b00000000 ;
			15'h00004203 : data <= 8'b00000000 ;
			15'h00004204 : data <= 8'b00000000 ;
			15'h00004205 : data <= 8'b00000000 ;
			15'h00004206 : data <= 8'b00000000 ;
			15'h00004207 : data <= 8'b00000000 ;
			15'h00004208 : data <= 8'b00000000 ;
			15'h00004209 : data <= 8'b00000000 ;
			15'h0000420A : data <= 8'b00000000 ;
			15'h0000420B : data <= 8'b00000000 ;
			15'h0000420C : data <= 8'b00000000 ;
			15'h0000420D : data <= 8'b00000000 ;
			15'h0000420E : data <= 8'b00000000 ;
			15'h0000420F : data <= 8'b00000000 ;
			15'h00004210 : data <= 8'b00000000 ;
			15'h00004211 : data <= 8'b00000000 ;
			15'h00004212 : data <= 8'b00000000 ;
			15'h00004213 : data <= 8'b00000000 ;
			15'h00004214 : data <= 8'b00000000 ;
			15'h00004215 : data <= 8'b00000000 ;
			15'h00004216 : data <= 8'b00000000 ;
			15'h00004217 : data <= 8'b00000000 ;
			15'h00004218 : data <= 8'b00000000 ;
			15'h00004219 : data <= 8'b00000000 ;
			15'h0000421A : data <= 8'b00000000 ;
			15'h0000421B : data <= 8'b00000000 ;
			15'h0000421C : data <= 8'b00000000 ;
			15'h0000421D : data <= 8'b00000000 ;
			15'h0000421E : data <= 8'b00000000 ;
			15'h0000421F : data <= 8'b00000000 ;
			15'h00004220 : data <= 8'b00000000 ;
			15'h00004221 : data <= 8'b00000000 ;
			15'h00004222 : data <= 8'b00000000 ;
			15'h00004223 : data <= 8'b00000000 ;
			15'h00004224 : data <= 8'b00000000 ;
			15'h00004225 : data <= 8'b00000000 ;
			15'h00004226 : data <= 8'b00000000 ;
			15'h00004227 : data <= 8'b00000000 ;
			15'h00004228 : data <= 8'b00000000 ;
			15'h00004229 : data <= 8'b00000000 ;
			15'h0000422A : data <= 8'b00000000 ;
			15'h0000422B : data <= 8'b00000000 ;
			15'h0000422C : data <= 8'b00000000 ;
			15'h0000422D : data <= 8'b00000000 ;
			15'h0000422E : data <= 8'b00000000 ;
			15'h0000422F : data <= 8'b00000000 ;
			15'h00004230 : data <= 8'b00000000 ;
			15'h00004231 : data <= 8'b00000000 ;
			15'h00004232 : data <= 8'b00000000 ;
			15'h00004233 : data <= 8'b00000000 ;
			15'h00004234 : data <= 8'b00000000 ;
			15'h00004235 : data <= 8'b00000000 ;
			15'h00004236 : data <= 8'b00000000 ;
			15'h00004237 : data <= 8'b00000000 ;
			15'h00004238 : data <= 8'b00000000 ;
			15'h00004239 : data <= 8'b00000000 ;
			15'h0000423A : data <= 8'b00000000 ;
			15'h0000423B : data <= 8'b00000000 ;
			15'h0000423C : data <= 8'b00000000 ;
			15'h0000423D : data <= 8'b00000000 ;
			15'h0000423E : data <= 8'b00000000 ;
			15'h0000423F : data <= 8'b00000000 ;
			15'h00004240 : data <= 8'b00000000 ;
			15'h00004241 : data <= 8'b00000000 ;
			15'h00004242 : data <= 8'b00000000 ;
			15'h00004243 : data <= 8'b00000000 ;
			15'h00004244 : data <= 8'b00000000 ;
			15'h00004245 : data <= 8'b00000000 ;
			15'h00004246 : data <= 8'b00000000 ;
			15'h00004247 : data <= 8'b00000000 ;
			15'h00004248 : data <= 8'b00000000 ;
			15'h00004249 : data <= 8'b00000000 ;
			15'h0000424A : data <= 8'b00000000 ;
			15'h0000424B : data <= 8'b00000000 ;
			15'h0000424C : data <= 8'b00000000 ;
			15'h0000424D : data <= 8'b00000000 ;
			15'h0000424E : data <= 8'b00000000 ;
			15'h0000424F : data <= 8'b00000000 ;
			15'h00004250 : data <= 8'b00000000 ;
			15'h00004251 : data <= 8'b00000000 ;
			15'h00004252 : data <= 8'b00000000 ;
			15'h00004253 : data <= 8'b00000000 ;
			15'h00004254 : data <= 8'b00000000 ;
			15'h00004255 : data <= 8'b00000000 ;
			15'h00004256 : data <= 8'b00000000 ;
			15'h00004257 : data <= 8'b00000000 ;
			15'h00004258 : data <= 8'b00000000 ;
			15'h00004259 : data <= 8'b00000000 ;
			15'h0000425A : data <= 8'b00000000 ;
			15'h0000425B : data <= 8'b00000000 ;
			15'h0000425C : data <= 8'b00000000 ;
			15'h0000425D : data <= 8'b00000000 ;
			15'h0000425E : data <= 8'b00000000 ;
			15'h0000425F : data <= 8'b00000000 ;
			15'h00004260 : data <= 8'b00000000 ;
			15'h00004261 : data <= 8'b00000000 ;
			15'h00004262 : data <= 8'b00000000 ;
			15'h00004263 : data <= 8'b00000000 ;
			15'h00004264 : data <= 8'b00000000 ;
			15'h00004265 : data <= 8'b00000000 ;
			15'h00004266 : data <= 8'b00000000 ;
			15'h00004267 : data <= 8'b00000000 ;
			15'h00004268 : data <= 8'b00000000 ;
			15'h00004269 : data <= 8'b00000000 ;
			15'h0000426A : data <= 8'b00000000 ;
			15'h0000426B : data <= 8'b00000000 ;
			15'h0000426C : data <= 8'b00000000 ;
			15'h0000426D : data <= 8'b00000000 ;
			15'h0000426E : data <= 8'b00000000 ;
			15'h0000426F : data <= 8'b00000000 ;
			15'h00004270 : data <= 8'b00000000 ;
			15'h00004271 : data <= 8'b00000000 ;
			15'h00004272 : data <= 8'b00000000 ;
			15'h00004273 : data <= 8'b00000000 ;
			15'h00004274 : data <= 8'b00000000 ;
			15'h00004275 : data <= 8'b00000000 ;
			15'h00004276 : data <= 8'b00000000 ;
			15'h00004277 : data <= 8'b00000000 ;
			15'h00004278 : data <= 8'b00000000 ;
			15'h00004279 : data <= 8'b00000000 ;
			15'h0000427A : data <= 8'b00000000 ;
			15'h0000427B : data <= 8'b00000000 ;
			15'h0000427C : data <= 8'b00000000 ;
			15'h0000427D : data <= 8'b00000000 ;
			15'h0000427E : data <= 8'b00000000 ;
			15'h0000427F : data <= 8'b00000000 ;
			15'h00004280 : data <= 8'b00000000 ;
			15'h00004281 : data <= 8'b00000000 ;
			15'h00004282 : data <= 8'b00000000 ;
			15'h00004283 : data <= 8'b00000000 ;
			15'h00004284 : data <= 8'b00000000 ;
			15'h00004285 : data <= 8'b00000000 ;
			15'h00004286 : data <= 8'b00000000 ;
			15'h00004287 : data <= 8'b00000000 ;
			15'h00004288 : data <= 8'b00000000 ;
			15'h00004289 : data <= 8'b00000000 ;
			15'h0000428A : data <= 8'b00000000 ;
			15'h0000428B : data <= 8'b00000000 ;
			15'h0000428C : data <= 8'b00000000 ;
			15'h0000428D : data <= 8'b00000000 ;
			15'h0000428E : data <= 8'b00000000 ;
			15'h0000428F : data <= 8'b00000000 ;
			15'h00004290 : data <= 8'b00000000 ;
			15'h00004291 : data <= 8'b00000000 ;
			15'h00004292 : data <= 8'b00000000 ;
			15'h00004293 : data <= 8'b00000000 ;
			15'h00004294 : data <= 8'b00000000 ;
			15'h00004295 : data <= 8'b00000000 ;
			15'h00004296 : data <= 8'b00000000 ;
			15'h00004297 : data <= 8'b00000000 ;
			15'h00004298 : data <= 8'b00000000 ;
			15'h00004299 : data <= 8'b00000000 ;
			15'h0000429A : data <= 8'b00000000 ;
			15'h0000429B : data <= 8'b00000000 ;
			15'h0000429C : data <= 8'b00000000 ;
			15'h0000429D : data <= 8'b00000000 ;
			15'h0000429E : data <= 8'b00000000 ;
			15'h0000429F : data <= 8'b00000000 ;
			15'h000042A0 : data <= 8'b00000000 ;
			15'h000042A1 : data <= 8'b00000000 ;
			15'h000042A2 : data <= 8'b00000000 ;
			15'h000042A3 : data <= 8'b00000000 ;
			15'h000042A4 : data <= 8'b00000000 ;
			15'h000042A5 : data <= 8'b00000000 ;
			15'h000042A6 : data <= 8'b00000000 ;
			15'h000042A7 : data <= 8'b00000000 ;
			15'h000042A8 : data <= 8'b00000000 ;
			15'h000042A9 : data <= 8'b00000000 ;
			15'h000042AA : data <= 8'b00000000 ;
			15'h000042AB : data <= 8'b00000000 ;
			15'h000042AC : data <= 8'b00000000 ;
			15'h000042AD : data <= 8'b00000000 ;
			15'h000042AE : data <= 8'b00000000 ;
			15'h000042AF : data <= 8'b00000000 ;
			15'h000042B0 : data <= 8'b00000000 ;
			15'h000042B1 : data <= 8'b00000000 ;
			15'h000042B2 : data <= 8'b00000000 ;
			15'h000042B3 : data <= 8'b00000000 ;
			15'h000042B4 : data <= 8'b00000000 ;
			15'h000042B5 : data <= 8'b00000000 ;
			15'h000042B6 : data <= 8'b00000000 ;
			15'h000042B7 : data <= 8'b00000000 ;
			15'h000042B8 : data <= 8'b00000000 ;
			15'h000042B9 : data <= 8'b00000000 ;
			15'h000042BA : data <= 8'b00000000 ;
			15'h000042BB : data <= 8'b00000000 ;
			15'h000042BC : data <= 8'b00000000 ;
			15'h000042BD : data <= 8'b00000000 ;
			15'h000042BE : data <= 8'b00000000 ;
			15'h000042BF : data <= 8'b00000000 ;
			15'h000042C0 : data <= 8'b00000000 ;
			15'h000042C1 : data <= 8'b00000000 ;
			15'h000042C2 : data <= 8'b00000000 ;
			15'h000042C3 : data <= 8'b00000000 ;
			15'h000042C4 : data <= 8'b00000000 ;
			15'h000042C5 : data <= 8'b00000000 ;
			15'h000042C6 : data <= 8'b00000000 ;
			15'h000042C7 : data <= 8'b00000000 ;
			15'h000042C8 : data <= 8'b00000000 ;
			15'h000042C9 : data <= 8'b00000000 ;
			15'h000042CA : data <= 8'b00000000 ;
			15'h000042CB : data <= 8'b00000000 ;
			15'h000042CC : data <= 8'b00000000 ;
			15'h000042CD : data <= 8'b00000000 ;
			15'h000042CE : data <= 8'b00000000 ;
			15'h000042CF : data <= 8'b00000000 ;
			15'h000042D0 : data <= 8'b00000000 ;
			15'h000042D1 : data <= 8'b00000000 ;
			15'h000042D2 : data <= 8'b00000000 ;
			15'h000042D3 : data <= 8'b00000000 ;
			15'h000042D4 : data <= 8'b00000000 ;
			15'h000042D5 : data <= 8'b00000000 ;
			15'h000042D6 : data <= 8'b00000000 ;
			15'h000042D7 : data <= 8'b00000000 ;
			15'h000042D8 : data <= 8'b00000000 ;
			15'h000042D9 : data <= 8'b00000000 ;
			15'h000042DA : data <= 8'b00000000 ;
			15'h000042DB : data <= 8'b00000000 ;
			15'h000042DC : data <= 8'b00000000 ;
			15'h000042DD : data <= 8'b00000000 ;
			15'h000042DE : data <= 8'b00000000 ;
			15'h000042DF : data <= 8'b00000000 ;
			15'h000042E0 : data <= 8'b00000000 ;
			15'h000042E1 : data <= 8'b00000000 ;
			15'h000042E2 : data <= 8'b00000000 ;
			15'h000042E3 : data <= 8'b00000000 ;
			15'h000042E4 : data <= 8'b00000000 ;
			15'h000042E5 : data <= 8'b00000000 ;
			15'h000042E6 : data <= 8'b00000000 ;
			15'h000042E7 : data <= 8'b00000000 ;
			15'h000042E8 : data <= 8'b00000000 ;
			15'h000042E9 : data <= 8'b00000000 ;
			15'h000042EA : data <= 8'b00000000 ;
			15'h000042EB : data <= 8'b00000000 ;
			15'h000042EC : data <= 8'b00000000 ;
			15'h000042ED : data <= 8'b00000000 ;
			15'h000042EE : data <= 8'b00000000 ;
			15'h000042EF : data <= 8'b00000000 ;
			15'h000042F0 : data <= 8'b00000000 ;
			15'h000042F1 : data <= 8'b00000000 ;
			15'h000042F2 : data <= 8'b00000000 ;
			15'h000042F3 : data <= 8'b00000000 ;
			15'h000042F4 : data <= 8'b00000000 ;
			15'h000042F5 : data <= 8'b00000000 ;
			15'h000042F6 : data <= 8'b00000000 ;
			15'h000042F7 : data <= 8'b00000000 ;
			15'h000042F8 : data <= 8'b00000000 ;
			15'h000042F9 : data <= 8'b00000000 ;
			15'h000042FA : data <= 8'b00000000 ;
			15'h000042FB : data <= 8'b00000000 ;
			15'h000042FC : data <= 8'b00000000 ;
			15'h000042FD : data <= 8'b00000000 ;
			15'h000042FE : data <= 8'b00000000 ;
			15'h000042FF : data <= 8'b00000000 ;
			15'h00004300 : data <= 8'b00000000 ;
			15'h00004301 : data <= 8'b00000000 ;
			15'h00004302 : data <= 8'b00000000 ;
			15'h00004303 : data <= 8'b00000000 ;
			15'h00004304 : data <= 8'b00000000 ;
			15'h00004305 : data <= 8'b00000000 ;
			15'h00004306 : data <= 8'b00000000 ;
			15'h00004307 : data <= 8'b00000000 ;
			15'h00004308 : data <= 8'b00000000 ;
			15'h00004309 : data <= 8'b00000000 ;
			15'h0000430A : data <= 8'b00000000 ;
			15'h0000430B : data <= 8'b00000000 ;
			15'h0000430C : data <= 8'b00000000 ;
			15'h0000430D : data <= 8'b00000000 ;
			15'h0000430E : data <= 8'b00000000 ;
			15'h0000430F : data <= 8'b00000000 ;
			15'h00004310 : data <= 8'b00000000 ;
			15'h00004311 : data <= 8'b00000000 ;
			15'h00004312 : data <= 8'b00000000 ;
			15'h00004313 : data <= 8'b00000000 ;
			15'h00004314 : data <= 8'b00000000 ;
			15'h00004315 : data <= 8'b00000000 ;
			15'h00004316 : data <= 8'b00000000 ;
			15'h00004317 : data <= 8'b00000000 ;
			15'h00004318 : data <= 8'b00000000 ;
			15'h00004319 : data <= 8'b00000000 ;
			15'h0000431A : data <= 8'b00000000 ;
			15'h0000431B : data <= 8'b00000000 ;
			15'h0000431C : data <= 8'b00000000 ;
			15'h0000431D : data <= 8'b00000000 ;
			15'h0000431E : data <= 8'b00000000 ;
			15'h0000431F : data <= 8'b00000000 ;
			15'h00004320 : data <= 8'b00000000 ;
			15'h00004321 : data <= 8'b00000000 ;
			15'h00004322 : data <= 8'b00000000 ;
			15'h00004323 : data <= 8'b00000000 ;
			15'h00004324 : data <= 8'b00000000 ;
			15'h00004325 : data <= 8'b00000000 ;
			15'h00004326 : data <= 8'b00000000 ;
			15'h00004327 : data <= 8'b00000000 ;
			15'h00004328 : data <= 8'b00000000 ;
			15'h00004329 : data <= 8'b00000000 ;
			15'h0000432A : data <= 8'b00000000 ;
			15'h0000432B : data <= 8'b00000000 ;
			15'h0000432C : data <= 8'b00000000 ;
			15'h0000432D : data <= 8'b00000000 ;
			15'h0000432E : data <= 8'b00000000 ;
			15'h0000432F : data <= 8'b00000000 ;
			15'h00004330 : data <= 8'b00000000 ;
			15'h00004331 : data <= 8'b00000000 ;
			15'h00004332 : data <= 8'b00000000 ;
			15'h00004333 : data <= 8'b00000000 ;
			15'h00004334 : data <= 8'b00000000 ;
			15'h00004335 : data <= 8'b00000000 ;
			15'h00004336 : data <= 8'b00000000 ;
			15'h00004337 : data <= 8'b00000000 ;
			15'h00004338 : data <= 8'b00000000 ;
			15'h00004339 : data <= 8'b00000000 ;
			15'h0000433A : data <= 8'b00000000 ;
			15'h0000433B : data <= 8'b00000000 ;
			15'h0000433C : data <= 8'b00000000 ;
			15'h0000433D : data <= 8'b00000000 ;
			15'h0000433E : data <= 8'b00000000 ;
			15'h0000433F : data <= 8'b00000000 ;
			15'h00004340 : data <= 8'b00000000 ;
			15'h00004341 : data <= 8'b00000000 ;
			15'h00004342 : data <= 8'b00000000 ;
			15'h00004343 : data <= 8'b00000000 ;
			15'h00004344 : data <= 8'b00000000 ;
			15'h00004345 : data <= 8'b00000000 ;
			15'h00004346 : data <= 8'b00000000 ;
			15'h00004347 : data <= 8'b00000000 ;
			15'h00004348 : data <= 8'b00000000 ;
			15'h00004349 : data <= 8'b00000000 ;
			15'h0000434A : data <= 8'b00000000 ;
			15'h0000434B : data <= 8'b00000000 ;
			15'h0000434C : data <= 8'b00000000 ;
			15'h0000434D : data <= 8'b00000000 ;
			15'h0000434E : data <= 8'b00000000 ;
			15'h0000434F : data <= 8'b00000000 ;
			15'h00004350 : data <= 8'b00000000 ;
			15'h00004351 : data <= 8'b00000000 ;
			15'h00004352 : data <= 8'b00000000 ;
			15'h00004353 : data <= 8'b00000000 ;
			15'h00004354 : data <= 8'b00000000 ;
			15'h00004355 : data <= 8'b00000000 ;
			15'h00004356 : data <= 8'b00000000 ;
			15'h00004357 : data <= 8'b00000000 ;
			15'h00004358 : data <= 8'b00000000 ;
			15'h00004359 : data <= 8'b00000000 ;
			15'h0000435A : data <= 8'b00000000 ;
			15'h0000435B : data <= 8'b00000000 ;
			15'h0000435C : data <= 8'b00000000 ;
			15'h0000435D : data <= 8'b00000000 ;
			15'h0000435E : data <= 8'b00000000 ;
			15'h0000435F : data <= 8'b00000000 ;
			15'h00004360 : data <= 8'b00000000 ;
			15'h00004361 : data <= 8'b00000000 ;
			15'h00004362 : data <= 8'b00000000 ;
			15'h00004363 : data <= 8'b00000000 ;
			15'h00004364 : data <= 8'b00000000 ;
			15'h00004365 : data <= 8'b00000000 ;
			15'h00004366 : data <= 8'b00000000 ;
			15'h00004367 : data <= 8'b00000000 ;
			15'h00004368 : data <= 8'b00000000 ;
			15'h00004369 : data <= 8'b00000000 ;
			15'h0000436A : data <= 8'b00000000 ;
			15'h0000436B : data <= 8'b00000000 ;
			15'h0000436C : data <= 8'b00000000 ;
			15'h0000436D : data <= 8'b00000000 ;
			15'h0000436E : data <= 8'b00000000 ;
			15'h0000436F : data <= 8'b00000000 ;
			15'h00004370 : data <= 8'b00000000 ;
			15'h00004371 : data <= 8'b00000000 ;
			15'h00004372 : data <= 8'b00000000 ;
			15'h00004373 : data <= 8'b00000000 ;
			15'h00004374 : data <= 8'b00000000 ;
			15'h00004375 : data <= 8'b00000000 ;
			15'h00004376 : data <= 8'b00000000 ;
			15'h00004377 : data <= 8'b00000000 ;
			15'h00004378 : data <= 8'b00000000 ;
			15'h00004379 : data <= 8'b00000000 ;
			15'h0000437A : data <= 8'b00000000 ;
			15'h0000437B : data <= 8'b00000000 ;
			15'h0000437C : data <= 8'b00000000 ;
			15'h0000437D : data <= 8'b00000000 ;
			15'h0000437E : data <= 8'b00000000 ;
			15'h0000437F : data <= 8'b00000000 ;
			15'h00004380 : data <= 8'b00000000 ;
			15'h00004381 : data <= 8'b00000000 ;
			15'h00004382 : data <= 8'b00000000 ;
			15'h00004383 : data <= 8'b00000000 ;
			15'h00004384 : data <= 8'b00000000 ;
			15'h00004385 : data <= 8'b00000000 ;
			15'h00004386 : data <= 8'b00000000 ;
			15'h00004387 : data <= 8'b00000000 ;
			15'h00004388 : data <= 8'b00000000 ;
			15'h00004389 : data <= 8'b00000000 ;
			15'h0000438A : data <= 8'b00000000 ;
			15'h0000438B : data <= 8'b00000000 ;
			15'h0000438C : data <= 8'b00000000 ;
			15'h0000438D : data <= 8'b00000000 ;
			15'h0000438E : data <= 8'b00000000 ;
			15'h0000438F : data <= 8'b00000000 ;
			15'h00004390 : data <= 8'b00000000 ;
			15'h00004391 : data <= 8'b00000000 ;
			15'h00004392 : data <= 8'b00000000 ;
			15'h00004393 : data <= 8'b00000000 ;
			15'h00004394 : data <= 8'b00000000 ;
			15'h00004395 : data <= 8'b00000000 ;
			15'h00004396 : data <= 8'b00000000 ;
			15'h00004397 : data <= 8'b00000000 ;
			15'h00004398 : data <= 8'b00000000 ;
			15'h00004399 : data <= 8'b00000000 ;
			15'h0000439A : data <= 8'b00000000 ;
			15'h0000439B : data <= 8'b00000000 ;
			15'h0000439C : data <= 8'b00000000 ;
			15'h0000439D : data <= 8'b00000000 ;
			15'h0000439E : data <= 8'b00000000 ;
			15'h0000439F : data <= 8'b00000000 ;
			15'h000043A0 : data <= 8'b00000000 ;
			15'h000043A1 : data <= 8'b00000000 ;
			15'h000043A2 : data <= 8'b00000000 ;
			15'h000043A3 : data <= 8'b00000000 ;
			15'h000043A4 : data <= 8'b00000000 ;
			15'h000043A5 : data <= 8'b00000000 ;
			15'h000043A6 : data <= 8'b00000000 ;
			15'h000043A7 : data <= 8'b00000000 ;
			15'h000043A8 : data <= 8'b00000000 ;
			15'h000043A9 : data <= 8'b00000000 ;
			15'h000043AA : data <= 8'b00000000 ;
			15'h000043AB : data <= 8'b00000000 ;
			15'h000043AC : data <= 8'b00000000 ;
			15'h000043AD : data <= 8'b00000000 ;
			15'h000043AE : data <= 8'b00000000 ;
			15'h000043AF : data <= 8'b00000000 ;
			15'h000043B0 : data <= 8'b00000000 ;
			15'h000043B1 : data <= 8'b00000000 ;
			15'h000043B2 : data <= 8'b00000000 ;
			15'h000043B3 : data <= 8'b00000000 ;
			15'h000043B4 : data <= 8'b00000000 ;
			15'h000043B5 : data <= 8'b00000000 ;
			15'h000043B6 : data <= 8'b00000000 ;
			15'h000043B7 : data <= 8'b00000000 ;
			15'h000043B8 : data <= 8'b00000000 ;
			15'h000043B9 : data <= 8'b00000000 ;
			15'h000043BA : data <= 8'b00000000 ;
			15'h000043BB : data <= 8'b00000000 ;
			15'h000043BC : data <= 8'b00000000 ;
			15'h000043BD : data <= 8'b00000000 ;
			15'h000043BE : data <= 8'b00000000 ;
			15'h000043BF : data <= 8'b00000000 ;
			15'h000043C0 : data <= 8'b00000000 ;
			15'h000043C1 : data <= 8'b00000000 ;
			15'h000043C2 : data <= 8'b00000000 ;
			15'h000043C3 : data <= 8'b00000000 ;
			15'h000043C4 : data <= 8'b00000000 ;
			15'h000043C5 : data <= 8'b00000000 ;
			15'h000043C6 : data <= 8'b00000000 ;
			15'h000043C7 : data <= 8'b00000000 ;
			15'h000043C8 : data <= 8'b00000000 ;
			15'h000043C9 : data <= 8'b00000000 ;
			15'h000043CA : data <= 8'b00000000 ;
			15'h000043CB : data <= 8'b00000000 ;
			15'h000043CC : data <= 8'b00000000 ;
			15'h000043CD : data <= 8'b00000000 ;
			15'h000043CE : data <= 8'b00000000 ;
			15'h000043CF : data <= 8'b00000000 ;
			15'h000043D0 : data <= 8'b00000000 ;
			15'h000043D1 : data <= 8'b00000000 ;
			15'h000043D2 : data <= 8'b00000000 ;
			15'h000043D3 : data <= 8'b00000000 ;
			15'h000043D4 : data <= 8'b00000000 ;
			15'h000043D5 : data <= 8'b00000000 ;
			15'h000043D6 : data <= 8'b00000000 ;
			15'h000043D7 : data <= 8'b00000000 ;
			15'h000043D8 : data <= 8'b00000000 ;
			15'h000043D9 : data <= 8'b00000000 ;
			15'h000043DA : data <= 8'b00000000 ;
			15'h000043DB : data <= 8'b00000000 ;
			15'h000043DC : data <= 8'b00000000 ;
			15'h000043DD : data <= 8'b00000000 ;
			15'h000043DE : data <= 8'b00000000 ;
			15'h000043DF : data <= 8'b00000000 ;
			15'h000043E0 : data <= 8'b00000000 ;
			15'h000043E1 : data <= 8'b00000000 ;
			15'h000043E2 : data <= 8'b00000000 ;
			15'h000043E3 : data <= 8'b00000000 ;
			15'h000043E4 : data <= 8'b00000000 ;
			15'h000043E5 : data <= 8'b00000000 ;
			15'h000043E6 : data <= 8'b00000000 ;
			15'h000043E7 : data <= 8'b00000000 ;
			15'h000043E8 : data <= 8'b00000000 ;
			15'h000043E9 : data <= 8'b00000000 ;
			15'h000043EA : data <= 8'b00000000 ;
			15'h000043EB : data <= 8'b00000000 ;
			15'h000043EC : data <= 8'b00000000 ;
			15'h000043ED : data <= 8'b00000000 ;
			15'h000043EE : data <= 8'b00000000 ;
			15'h000043EF : data <= 8'b00000000 ;
			15'h000043F0 : data <= 8'b00000000 ;
			15'h000043F1 : data <= 8'b00000000 ;
			15'h000043F2 : data <= 8'b00000000 ;
			15'h000043F3 : data <= 8'b00000000 ;
			15'h000043F4 : data <= 8'b00000000 ;
			15'h000043F5 : data <= 8'b00000000 ;
			15'h000043F6 : data <= 8'b00000000 ;
			15'h000043F7 : data <= 8'b00000000 ;
			15'h000043F8 : data <= 8'b00000000 ;
			15'h000043F9 : data <= 8'b00000000 ;
			15'h000043FA : data <= 8'b00000000 ;
			15'h000043FB : data <= 8'b00000000 ;
			15'h000043FC : data <= 8'b00000000 ;
			15'h000043FD : data <= 8'b00000000 ;
			15'h000043FE : data <= 8'b00000000 ;
			15'h000043FF : data <= 8'b00000000 ;
			15'h00004400 : data <= 8'b00000000 ;
			15'h00004401 : data <= 8'b00000000 ;
			15'h00004402 : data <= 8'b00000000 ;
			15'h00004403 : data <= 8'b00000000 ;
			15'h00004404 : data <= 8'b00000000 ;
			15'h00004405 : data <= 8'b00000000 ;
			15'h00004406 : data <= 8'b00000000 ;
			15'h00004407 : data <= 8'b00000000 ;
			15'h00004408 : data <= 8'b00000000 ;
			15'h00004409 : data <= 8'b00000000 ;
			15'h0000440A : data <= 8'b00000000 ;
			15'h0000440B : data <= 8'b00000000 ;
			15'h0000440C : data <= 8'b00000000 ;
			15'h0000440D : data <= 8'b00000000 ;
			15'h0000440E : data <= 8'b00000000 ;
			15'h0000440F : data <= 8'b00000000 ;
			15'h00004410 : data <= 8'b00000000 ;
			15'h00004411 : data <= 8'b00000000 ;
			15'h00004412 : data <= 8'b00000000 ;
			15'h00004413 : data <= 8'b00000000 ;
			15'h00004414 : data <= 8'b00000000 ;
			15'h00004415 : data <= 8'b00000000 ;
			15'h00004416 : data <= 8'b00000000 ;
			15'h00004417 : data <= 8'b00000000 ;
			15'h00004418 : data <= 8'b00000000 ;
			15'h00004419 : data <= 8'b00000000 ;
			15'h0000441A : data <= 8'b00000000 ;
			15'h0000441B : data <= 8'b00000000 ;
			15'h0000441C : data <= 8'b00000000 ;
			15'h0000441D : data <= 8'b00000000 ;
			15'h0000441E : data <= 8'b00000000 ;
			15'h0000441F : data <= 8'b00000000 ;
			15'h00004420 : data <= 8'b00000000 ;
			15'h00004421 : data <= 8'b00000000 ;
			15'h00004422 : data <= 8'b00000000 ;
			15'h00004423 : data <= 8'b00000000 ;
			15'h00004424 : data <= 8'b00000000 ;
			15'h00004425 : data <= 8'b00000000 ;
			15'h00004426 : data <= 8'b00000000 ;
			15'h00004427 : data <= 8'b00000000 ;
			15'h00004428 : data <= 8'b00000000 ;
			15'h00004429 : data <= 8'b00000000 ;
			15'h0000442A : data <= 8'b00000000 ;
			15'h0000442B : data <= 8'b00000000 ;
			15'h0000442C : data <= 8'b00000000 ;
			15'h0000442D : data <= 8'b00000000 ;
			15'h0000442E : data <= 8'b00000000 ;
			15'h0000442F : data <= 8'b00000000 ;
			15'h00004430 : data <= 8'b00000000 ;
			15'h00004431 : data <= 8'b00000000 ;
			15'h00004432 : data <= 8'b00000000 ;
			15'h00004433 : data <= 8'b00000000 ;
			15'h00004434 : data <= 8'b00000000 ;
			15'h00004435 : data <= 8'b00000000 ;
			15'h00004436 : data <= 8'b00000000 ;
			15'h00004437 : data <= 8'b00000000 ;
			15'h00004438 : data <= 8'b00000000 ;
			15'h00004439 : data <= 8'b00000000 ;
			15'h0000443A : data <= 8'b00000000 ;
			15'h0000443B : data <= 8'b00000000 ;
			15'h0000443C : data <= 8'b00000000 ;
			15'h0000443D : data <= 8'b00000000 ;
			15'h0000443E : data <= 8'b00000000 ;
			15'h0000443F : data <= 8'b00000000 ;
			15'h00004440 : data <= 8'b00000000 ;
			15'h00004441 : data <= 8'b00000000 ;
			15'h00004442 : data <= 8'b00000000 ;
			15'h00004443 : data <= 8'b00000000 ;
			15'h00004444 : data <= 8'b00000000 ;
			15'h00004445 : data <= 8'b00000000 ;
			15'h00004446 : data <= 8'b00000000 ;
			15'h00004447 : data <= 8'b00000000 ;
			15'h00004448 : data <= 8'b00000000 ;
			15'h00004449 : data <= 8'b00000000 ;
			15'h0000444A : data <= 8'b00000000 ;
			15'h0000444B : data <= 8'b00000000 ;
			15'h0000444C : data <= 8'b00000000 ;
			15'h0000444D : data <= 8'b00000000 ;
			15'h0000444E : data <= 8'b00000000 ;
			15'h0000444F : data <= 8'b00000000 ;
			15'h00004450 : data <= 8'b00000000 ;
			15'h00004451 : data <= 8'b00000000 ;
			15'h00004452 : data <= 8'b00000000 ;
			15'h00004453 : data <= 8'b00000000 ;
			15'h00004454 : data <= 8'b00000000 ;
			15'h00004455 : data <= 8'b00000000 ;
			15'h00004456 : data <= 8'b00000000 ;
			15'h00004457 : data <= 8'b00000000 ;
			15'h00004458 : data <= 8'b00000000 ;
			15'h00004459 : data <= 8'b00000000 ;
			15'h0000445A : data <= 8'b00000000 ;
			15'h0000445B : data <= 8'b00000000 ;
			15'h0000445C : data <= 8'b00000000 ;
			15'h0000445D : data <= 8'b00000000 ;
			15'h0000445E : data <= 8'b00000000 ;
			15'h0000445F : data <= 8'b00000000 ;
			15'h00004460 : data <= 8'b00000000 ;
			15'h00004461 : data <= 8'b00000000 ;
			15'h00004462 : data <= 8'b00000000 ;
			15'h00004463 : data <= 8'b00000000 ;
			15'h00004464 : data <= 8'b00000000 ;
			15'h00004465 : data <= 8'b00000000 ;
			15'h00004466 : data <= 8'b00000000 ;
			15'h00004467 : data <= 8'b00000000 ;
			15'h00004468 : data <= 8'b00000000 ;
			15'h00004469 : data <= 8'b00000000 ;
			15'h0000446A : data <= 8'b00000000 ;
			15'h0000446B : data <= 8'b00000000 ;
			15'h0000446C : data <= 8'b00000000 ;
			15'h0000446D : data <= 8'b00000000 ;
			15'h0000446E : data <= 8'b00000000 ;
			15'h0000446F : data <= 8'b00000000 ;
			15'h00004470 : data <= 8'b00000000 ;
			15'h00004471 : data <= 8'b00000000 ;
			15'h00004472 : data <= 8'b00000000 ;
			15'h00004473 : data <= 8'b00000000 ;
			15'h00004474 : data <= 8'b00000000 ;
			15'h00004475 : data <= 8'b00000000 ;
			15'h00004476 : data <= 8'b00000000 ;
			15'h00004477 : data <= 8'b00000000 ;
			15'h00004478 : data <= 8'b00000000 ;
			15'h00004479 : data <= 8'b00000000 ;
			15'h0000447A : data <= 8'b00000000 ;
			15'h0000447B : data <= 8'b00000000 ;
			15'h0000447C : data <= 8'b00000000 ;
			15'h0000447D : data <= 8'b00000000 ;
			15'h0000447E : data <= 8'b00000000 ;
			15'h0000447F : data <= 8'b00000000 ;
			15'h00004480 : data <= 8'b00000000 ;
			15'h00004481 : data <= 8'b00000000 ;
			15'h00004482 : data <= 8'b00000000 ;
			15'h00004483 : data <= 8'b00000000 ;
			15'h00004484 : data <= 8'b00000000 ;
			15'h00004485 : data <= 8'b00000000 ;
			15'h00004486 : data <= 8'b00000000 ;
			15'h00004487 : data <= 8'b00000000 ;
			15'h00004488 : data <= 8'b00000000 ;
			15'h00004489 : data <= 8'b00000000 ;
			15'h0000448A : data <= 8'b00000000 ;
			15'h0000448B : data <= 8'b00000000 ;
			15'h0000448C : data <= 8'b00000000 ;
			15'h0000448D : data <= 8'b00000000 ;
			15'h0000448E : data <= 8'b00000000 ;
			15'h0000448F : data <= 8'b00000000 ;
			15'h00004490 : data <= 8'b00000000 ;
			15'h00004491 : data <= 8'b00000000 ;
			15'h00004492 : data <= 8'b00000000 ;
			15'h00004493 : data <= 8'b00000000 ;
			15'h00004494 : data <= 8'b00000000 ;
			15'h00004495 : data <= 8'b00000000 ;
			15'h00004496 : data <= 8'b00000000 ;
			15'h00004497 : data <= 8'b00000000 ;
			15'h00004498 : data <= 8'b00000000 ;
			15'h00004499 : data <= 8'b00000000 ;
			15'h0000449A : data <= 8'b00000000 ;
			15'h0000449B : data <= 8'b00000000 ;
			15'h0000449C : data <= 8'b00000000 ;
			15'h0000449D : data <= 8'b00000000 ;
			15'h0000449E : data <= 8'b00000000 ;
			15'h0000449F : data <= 8'b00000000 ;
			15'h000044A0 : data <= 8'b00000000 ;
			15'h000044A1 : data <= 8'b00000000 ;
			15'h000044A2 : data <= 8'b00000000 ;
			15'h000044A3 : data <= 8'b00000000 ;
			15'h000044A4 : data <= 8'b00000000 ;
			15'h000044A5 : data <= 8'b00000000 ;
			15'h000044A6 : data <= 8'b00000000 ;
			15'h000044A7 : data <= 8'b00000000 ;
			15'h000044A8 : data <= 8'b00000000 ;
			15'h000044A9 : data <= 8'b00000000 ;
			15'h000044AA : data <= 8'b00000000 ;
			15'h000044AB : data <= 8'b00000000 ;
			15'h000044AC : data <= 8'b00000000 ;
			15'h000044AD : data <= 8'b00000000 ;
			15'h000044AE : data <= 8'b00000000 ;
			15'h000044AF : data <= 8'b00000000 ;
			15'h000044B0 : data <= 8'b00000000 ;
			15'h000044B1 : data <= 8'b00000000 ;
			15'h000044B2 : data <= 8'b00000000 ;
			15'h000044B3 : data <= 8'b00000000 ;
			15'h000044B4 : data <= 8'b00000000 ;
			15'h000044B5 : data <= 8'b00000000 ;
			15'h000044B6 : data <= 8'b00000000 ;
			15'h000044B7 : data <= 8'b00000000 ;
			15'h000044B8 : data <= 8'b00000000 ;
			15'h000044B9 : data <= 8'b00000000 ;
			15'h000044BA : data <= 8'b00000000 ;
			15'h000044BB : data <= 8'b00000000 ;
			15'h000044BC : data <= 8'b00000000 ;
			15'h000044BD : data <= 8'b00000000 ;
			15'h000044BE : data <= 8'b00000000 ;
			15'h000044BF : data <= 8'b00000000 ;
			15'h000044C0 : data <= 8'b00000000 ;
			15'h000044C1 : data <= 8'b00000000 ;
			15'h000044C2 : data <= 8'b00000000 ;
			15'h000044C3 : data <= 8'b00000000 ;
			15'h000044C4 : data <= 8'b00000000 ;
			15'h000044C5 : data <= 8'b00000000 ;
			15'h000044C6 : data <= 8'b00000000 ;
			15'h000044C7 : data <= 8'b00000000 ;
			15'h000044C8 : data <= 8'b00000000 ;
			15'h000044C9 : data <= 8'b00000000 ;
			15'h000044CA : data <= 8'b00000000 ;
			15'h000044CB : data <= 8'b00000000 ;
			15'h000044CC : data <= 8'b00000000 ;
			15'h000044CD : data <= 8'b00000000 ;
			15'h000044CE : data <= 8'b00000000 ;
			15'h000044CF : data <= 8'b00000000 ;
			15'h000044D0 : data <= 8'b00000000 ;
			15'h000044D1 : data <= 8'b00000000 ;
			15'h000044D2 : data <= 8'b00000000 ;
			15'h000044D3 : data <= 8'b00000000 ;
			15'h000044D4 : data <= 8'b00000000 ;
			15'h000044D5 : data <= 8'b00000000 ;
			15'h000044D6 : data <= 8'b00000000 ;
			15'h000044D7 : data <= 8'b00000000 ;
			15'h000044D8 : data <= 8'b00000000 ;
			15'h000044D9 : data <= 8'b00000000 ;
			15'h000044DA : data <= 8'b00000000 ;
			15'h000044DB : data <= 8'b00000000 ;
			15'h000044DC : data <= 8'b00000000 ;
			15'h000044DD : data <= 8'b00000000 ;
			15'h000044DE : data <= 8'b00000000 ;
			15'h000044DF : data <= 8'b00000000 ;
			15'h000044E0 : data <= 8'b00000000 ;
			15'h000044E1 : data <= 8'b00000000 ;
			15'h000044E2 : data <= 8'b00000000 ;
			15'h000044E3 : data <= 8'b00000000 ;
			15'h000044E4 : data <= 8'b00000000 ;
			15'h000044E5 : data <= 8'b00000000 ;
			15'h000044E6 : data <= 8'b00000000 ;
			15'h000044E7 : data <= 8'b00000000 ;
			15'h000044E8 : data <= 8'b00000000 ;
			15'h000044E9 : data <= 8'b00000000 ;
			15'h000044EA : data <= 8'b00000000 ;
			15'h000044EB : data <= 8'b00000000 ;
			15'h000044EC : data <= 8'b00000000 ;
			15'h000044ED : data <= 8'b00000000 ;
			15'h000044EE : data <= 8'b00000000 ;
			15'h000044EF : data <= 8'b00000000 ;
			15'h000044F0 : data <= 8'b00000000 ;
			15'h000044F1 : data <= 8'b00000000 ;
			15'h000044F2 : data <= 8'b00000000 ;
			15'h000044F3 : data <= 8'b00000000 ;
			15'h000044F4 : data <= 8'b00000000 ;
			15'h000044F5 : data <= 8'b00000000 ;
			15'h000044F6 : data <= 8'b00000000 ;
			15'h000044F7 : data <= 8'b00000000 ;
			15'h000044F8 : data <= 8'b00000000 ;
			15'h000044F9 : data <= 8'b00000000 ;
			15'h000044FA : data <= 8'b00000000 ;
			15'h000044FB : data <= 8'b00000000 ;
			15'h000044FC : data <= 8'b00000000 ;
			15'h000044FD : data <= 8'b00000000 ;
			15'h000044FE : data <= 8'b00000000 ;
			15'h000044FF : data <= 8'b00000000 ;
			15'h00004500 : data <= 8'b00000000 ;
			15'h00004501 : data <= 8'b00000000 ;
			15'h00004502 : data <= 8'b00000000 ;
			15'h00004503 : data <= 8'b00000000 ;
			15'h00004504 : data <= 8'b00000000 ;
			15'h00004505 : data <= 8'b00000000 ;
			15'h00004506 : data <= 8'b00000000 ;
			15'h00004507 : data <= 8'b00000000 ;
			15'h00004508 : data <= 8'b00000000 ;
			15'h00004509 : data <= 8'b00000000 ;
			15'h0000450A : data <= 8'b00000000 ;
			15'h0000450B : data <= 8'b00000000 ;
			15'h0000450C : data <= 8'b00000000 ;
			15'h0000450D : data <= 8'b00000000 ;
			15'h0000450E : data <= 8'b00000000 ;
			15'h0000450F : data <= 8'b00000000 ;
			15'h00004510 : data <= 8'b00000000 ;
			15'h00004511 : data <= 8'b00000000 ;
			15'h00004512 : data <= 8'b00000000 ;
			15'h00004513 : data <= 8'b00000000 ;
			15'h00004514 : data <= 8'b00000000 ;
			15'h00004515 : data <= 8'b00000000 ;
			15'h00004516 : data <= 8'b00000000 ;
			15'h00004517 : data <= 8'b00000000 ;
			15'h00004518 : data <= 8'b00000000 ;
			15'h00004519 : data <= 8'b00000000 ;
			15'h0000451A : data <= 8'b00000000 ;
			15'h0000451B : data <= 8'b00000000 ;
			15'h0000451C : data <= 8'b00000000 ;
			15'h0000451D : data <= 8'b00000000 ;
			15'h0000451E : data <= 8'b00000000 ;
			15'h0000451F : data <= 8'b00000000 ;
			15'h00004520 : data <= 8'b00000000 ;
			15'h00004521 : data <= 8'b00000000 ;
			15'h00004522 : data <= 8'b00000000 ;
			15'h00004523 : data <= 8'b00000000 ;
			15'h00004524 : data <= 8'b00000000 ;
			15'h00004525 : data <= 8'b00000000 ;
			15'h00004526 : data <= 8'b00000000 ;
			15'h00004527 : data <= 8'b00000000 ;
			15'h00004528 : data <= 8'b00000000 ;
			15'h00004529 : data <= 8'b00000000 ;
			15'h0000452A : data <= 8'b00000000 ;
			15'h0000452B : data <= 8'b00000000 ;
			15'h0000452C : data <= 8'b00000000 ;
			15'h0000452D : data <= 8'b00000000 ;
			15'h0000452E : data <= 8'b00000000 ;
			15'h0000452F : data <= 8'b00000000 ;
			15'h00004530 : data <= 8'b00000000 ;
			15'h00004531 : data <= 8'b00000000 ;
			15'h00004532 : data <= 8'b00000000 ;
			15'h00004533 : data <= 8'b00000000 ;
			15'h00004534 : data <= 8'b00000000 ;
			15'h00004535 : data <= 8'b00000000 ;
			15'h00004536 : data <= 8'b00000000 ;
			15'h00004537 : data <= 8'b00000000 ;
			15'h00004538 : data <= 8'b00000000 ;
			15'h00004539 : data <= 8'b00000000 ;
			15'h0000453A : data <= 8'b00000000 ;
			15'h0000453B : data <= 8'b00000000 ;
			15'h0000453C : data <= 8'b00000000 ;
			15'h0000453D : data <= 8'b00000000 ;
			15'h0000453E : data <= 8'b00000000 ;
			15'h0000453F : data <= 8'b00000000 ;
			15'h00004540 : data <= 8'b00000000 ;
			15'h00004541 : data <= 8'b00000000 ;
			15'h00004542 : data <= 8'b00000000 ;
			15'h00004543 : data <= 8'b00000000 ;
			15'h00004544 : data <= 8'b00000000 ;
			15'h00004545 : data <= 8'b00000000 ;
			15'h00004546 : data <= 8'b00000000 ;
			15'h00004547 : data <= 8'b00000000 ;
			15'h00004548 : data <= 8'b00000000 ;
			15'h00004549 : data <= 8'b00000000 ;
			15'h0000454A : data <= 8'b00000000 ;
			15'h0000454B : data <= 8'b00000000 ;
			15'h0000454C : data <= 8'b00000000 ;
			15'h0000454D : data <= 8'b00000000 ;
			15'h0000454E : data <= 8'b00000000 ;
			15'h0000454F : data <= 8'b00000000 ;
			15'h00004550 : data <= 8'b00000000 ;
			15'h00004551 : data <= 8'b00000000 ;
			15'h00004552 : data <= 8'b00000000 ;
			15'h00004553 : data <= 8'b00000000 ;
			15'h00004554 : data <= 8'b00000000 ;
			15'h00004555 : data <= 8'b00000000 ;
			15'h00004556 : data <= 8'b00000000 ;
			15'h00004557 : data <= 8'b00000000 ;
			15'h00004558 : data <= 8'b00000000 ;
			15'h00004559 : data <= 8'b00000000 ;
			15'h0000455A : data <= 8'b00000000 ;
			15'h0000455B : data <= 8'b00000000 ;
			15'h0000455C : data <= 8'b00000000 ;
			15'h0000455D : data <= 8'b00000000 ;
			15'h0000455E : data <= 8'b00000000 ;
			15'h0000455F : data <= 8'b00000000 ;
			15'h00004560 : data <= 8'b00000000 ;
			15'h00004561 : data <= 8'b00000000 ;
			15'h00004562 : data <= 8'b00000000 ;
			15'h00004563 : data <= 8'b00000000 ;
			15'h00004564 : data <= 8'b00000000 ;
			15'h00004565 : data <= 8'b00000000 ;
			15'h00004566 : data <= 8'b00000000 ;
			15'h00004567 : data <= 8'b00000000 ;
			15'h00004568 : data <= 8'b00000000 ;
			15'h00004569 : data <= 8'b00000000 ;
			15'h0000456A : data <= 8'b00000000 ;
			15'h0000456B : data <= 8'b00000000 ;
			15'h0000456C : data <= 8'b00000000 ;
			15'h0000456D : data <= 8'b00000000 ;
			15'h0000456E : data <= 8'b00000000 ;
			15'h0000456F : data <= 8'b00000000 ;
			15'h00004570 : data <= 8'b00000000 ;
			15'h00004571 : data <= 8'b00000000 ;
			15'h00004572 : data <= 8'b00000000 ;
			15'h00004573 : data <= 8'b00000000 ;
			15'h00004574 : data <= 8'b00000000 ;
			15'h00004575 : data <= 8'b00000000 ;
			15'h00004576 : data <= 8'b00000000 ;
			15'h00004577 : data <= 8'b00000000 ;
			15'h00004578 : data <= 8'b00000000 ;
			15'h00004579 : data <= 8'b00000000 ;
			15'h0000457A : data <= 8'b00000000 ;
			15'h0000457B : data <= 8'b00000000 ;
			15'h0000457C : data <= 8'b00000000 ;
			15'h0000457D : data <= 8'b00000000 ;
			15'h0000457E : data <= 8'b00000000 ;
			15'h0000457F : data <= 8'b00000000 ;
			15'h00004580 : data <= 8'b00000000 ;
			15'h00004581 : data <= 8'b00000000 ;
			15'h00004582 : data <= 8'b00000000 ;
			15'h00004583 : data <= 8'b00000000 ;
			15'h00004584 : data <= 8'b00000000 ;
			15'h00004585 : data <= 8'b00000000 ;
			15'h00004586 : data <= 8'b00000000 ;
			15'h00004587 : data <= 8'b00000000 ;
			15'h00004588 : data <= 8'b00000000 ;
			15'h00004589 : data <= 8'b00000000 ;
			15'h0000458A : data <= 8'b00000000 ;
			15'h0000458B : data <= 8'b00000000 ;
			15'h0000458C : data <= 8'b00000000 ;
			15'h0000458D : data <= 8'b00000000 ;
			15'h0000458E : data <= 8'b00000000 ;
			15'h0000458F : data <= 8'b00000000 ;
			15'h00004590 : data <= 8'b00000000 ;
			15'h00004591 : data <= 8'b00000000 ;
			15'h00004592 : data <= 8'b00000000 ;
			15'h00004593 : data <= 8'b00000000 ;
			15'h00004594 : data <= 8'b00000000 ;
			15'h00004595 : data <= 8'b00000000 ;
			15'h00004596 : data <= 8'b00000000 ;
			15'h00004597 : data <= 8'b00000000 ;
			15'h00004598 : data <= 8'b00000000 ;
			15'h00004599 : data <= 8'b00000000 ;
			15'h0000459A : data <= 8'b00000000 ;
			15'h0000459B : data <= 8'b00000000 ;
			15'h0000459C : data <= 8'b00000000 ;
			15'h0000459D : data <= 8'b00000000 ;
			15'h0000459E : data <= 8'b00000000 ;
			15'h0000459F : data <= 8'b00000000 ;
			15'h000045A0 : data <= 8'b00000000 ;
			15'h000045A1 : data <= 8'b00000000 ;
			15'h000045A2 : data <= 8'b00000000 ;
			15'h000045A3 : data <= 8'b00000000 ;
			15'h000045A4 : data <= 8'b00000000 ;
			15'h000045A5 : data <= 8'b00000000 ;
			15'h000045A6 : data <= 8'b00000000 ;
			15'h000045A7 : data <= 8'b00000000 ;
			15'h000045A8 : data <= 8'b00000000 ;
			15'h000045A9 : data <= 8'b00000000 ;
			15'h000045AA : data <= 8'b00000000 ;
			15'h000045AB : data <= 8'b00000000 ;
			15'h000045AC : data <= 8'b00000000 ;
			15'h000045AD : data <= 8'b00000000 ;
			15'h000045AE : data <= 8'b00000000 ;
			15'h000045AF : data <= 8'b00000000 ;
			15'h000045B0 : data <= 8'b00000000 ;
			15'h000045B1 : data <= 8'b00000000 ;
			15'h000045B2 : data <= 8'b00000000 ;
			15'h000045B3 : data <= 8'b00000000 ;
			15'h000045B4 : data <= 8'b00000000 ;
			15'h000045B5 : data <= 8'b00000000 ;
			15'h000045B6 : data <= 8'b00000000 ;
			15'h000045B7 : data <= 8'b00000000 ;
			15'h000045B8 : data <= 8'b00000000 ;
			15'h000045B9 : data <= 8'b00000000 ;
			15'h000045BA : data <= 8'b00000000 ;
			15'h000045BB : data <= 8'b00000000 ;
			15'h000045BC : data <= 8'b00000000 ;
			15'h000045BD : data <= 8'b00000000 ;
			15'h000045BE : data <= 8'b00000000 ;
			15'h000045BF : data <= 8'b00000000 ;
			15'h000045C0 : data <= 8'b00000000 ;
			15'h000045C1 : data <= 8'b00000000 ;
			15'h000045C2 : data <= 8'b00000000 ;
			15'h000045C3 : data <= 8'b00000000 ;
			15'h000045C4 : data <= 8'b00000000 ;
			15'h000045C5 : data <= 8'b00000000 ;
			15'h000045C6 : data <= 8'b00000000 ;
			15'h000045C7 : data <= 8'b00000000 ;
			15'h000045C8 : data <= 8'b00000000 ;
			15'h000045C9 : data <= 8'b00000000 ;
			15'h000045CA : data <= 8'b00000000 ;
			15'h000045CB : data <= 8'b00000000 ;
			15'h000045CC : data <= 8'b00000000 ;
			15'h000045CD : data <= 8'b00000000 ;
			15'h000045CE : data <= 8'b00000000 ;
			15'h000045CF : data <= 8'b00000000 ;
			15'h000045D0 : data <= 8'b00000000 ;
			15'h000045D1 : data <= 8'b00000000 ;
			15'h000045D2 : data <= 8'b00000000 ;
			15'h000045D3 : data <= 8'b00000000 ;
			15'h000045D4 : data <= 8'b00000000 ;
			15'h000045D5 : data <= 8'b00000000 ;
			15'h000045D6 : data <= 8'b00000000 ;
			15'h000045D7 : data <= 8'b00000000 ;
			15'h000045D8 : data <= 8'b00000000 ;
			15'h000045D9 : data <= 8'b00000000 ;
			15'h000045DA : data <= 8'b00000000 ;
			15'h000045DB : data <= 8'b00000000 ;
			15'h000045DC : data <= 8'b00000000 ;
			15'h000045DD : data <= 8'b00000000 ;
			15'h000045DE : data <= 8'b00000000 ;
			15'h000045DF : data <= 8'b00000000 ;
			15'h000045E0 : data <= 8'b00000000 ;
			15'h000045E1 : data <= 8'b00000000 ;
			15'h000045E2 : data <= 8'b00000000 ;
			15'h000045E3 : data <= 8'b00000000 ;
			15'h000045E4 : data <= 8'b00000000 ;
			15'h000045E5 : data <= 8'b00000000 ;
			15'h000045E6 : data <= 8'b00000000 ;
			15'h000045E7 : data <= 8'b00000000 ;
			15'h000045E8 : data <= 8'b00000000 ;
			15'h000045E9 : data <= 8'b00000000 ;
			15'h000045EA : data <= 8'b00000000 ;
			15'h000045EB : data <= 8'b00000000 ;
			15'h000045EC : data <= 8'b00000000 ;
			15'h000045ED : data <= 8'b00000000 ;
			15'h000045EE : data <= 8'b00000000 ;
			15'h000045EF : data <= 8'b00000000 ;
			15'h000045F0 : data <= 8'b00000000 ;
			15'h000045F1 : data <= 8'b00000000 ;
			15'h000045F2 : data <= 8'b00000000 ;
			15'h000045F3 : data <= 8'b00000000 ;
			15'h000045F4 : data <= 8'b00000000 ;
			15'h000045F5 : data <= 8'b00000000 ;
			15'h000045F6 : data <= 8'b00000000 ;
			15'h000045F7 : data <= 8'b00000000 ;
			15'h000045F8 : data <= 8'b00000000 ;
			15'h000045F9 : data <= 8'b00000000 ;
			15'h000045FA : data <= 8'b00000000 ;
			15'h000045FB : data <= 8'b00000000 ;
			15'h000045FC : data <= 8'b00000000 ;
			15'h000045FD : data <= 8'b00000000 ;
			15'h000045FE : data <= 8'b00000000 ;
			15'h000045FF : data <= 8'b00000000 ;
			15'h00004600 : data <= 8'b00000000 ;
			15'h00004601 : data <= 8'b00000000 ;
			15'h00004602 : data <= 8'b00000000 ;
			15'h00004603 : data <= 8'b00000000 ;
			15'h00004604 : data <= 8'b00000000 ;
			15'h00004605 : data <= 8'b00000000 ;
			15'h00004606 : data <= 8'b00000000 ;
			15'h00004607 : data <= 8'b00000000 ;
			15'h00004608 : data <= 8'b00000000 ;
			15'h00004609 : data <= 8'b00000000 ;
			15'h0000460A : data <= 8'b00000000 ;
			15'h0000460B : data <= 8'b00000000 ;
			15'h0000460C : data <= 8'b00000000 ;
			15'h0000460D : data <= 8'b00000000 ;
			15'h0000460E : data <= 8'b00000000 ;
			15'h0000460F : data <= 8'b00000000 ;
			15'h00004610 : data <= 8'b00000000 ;
			15'h00004611 : data <= 8'b00000000 ;
			15'h00004612 : data <= 8'b00000000 ;
			15'h00004613 : data <= 8'b00000000 ;
			15'h00004614 : data <= 8'b00000000 ;
			15'h00004615 : data <= 8'b00000000 ;
			15'h00004616 : data <= 8'b00000000 ;
			15'h00004617 : data <= 8'b00000000 ;
			15'h00004618 : data <= 8'b00000000 ;
			15'h00004619 : data <= 8'b00000000 ;
			15'h0000461A : data <= 8'b00000000 ;
			15'h0000461B : data <= 8'b00000000 ;
			15'h0000461C : data <= 8'b00000000 ;
			15'h0000461D : data <= 8'b00000000 ;
			15'h0000461E : data <= 8'b00000000 ;
			15'h0000461F : data <= 8'b00000000 ;
			15'h00004620 : data <= 8'b00000000 ;
			15'h00004621 : data <= 8'b00000000 ;
			15'h00004622 : data <= 8'b00000000 ;
			15'h00004623 : data <= 8'b00000000 ;
			15'h00004624 : data <= 8'b00000000 ;
			15'h00004625 : data <= 8'b00000000 ;
			15'h00004626 : data <= 8'b00000000 ;
			15'h00004627 : data <= 8'b00000000 ;
			15'h00004628 : data <= 8'b00000000 ;
			15'h00004629 : data <= 8'b00000000 ;
			15'h0000462A : data <= 8'b00000000 ;
			15'h0000462B : data <= 8'b00000000 ;
			15'h0000462C : data <= 8'b00000000 ;
			15'h0000462D : data <= 8'b00000000 ;
			15'h0000462E : data <= 8'b00000000 ;
			15'h0000462F : data <= 8'b00000000 ;
			15'h00004630 : data <= 8'b00000000 ;
			15'h00004631 : data <= 8'b00000000 ;
			15'h00004632 : data <= 8'b00000000 ;
			15'h00004633 : data <= 8'b00000000 ;
			15'h00004634 : data <= 8'b00000000 ;
			15'h00004635 : data <= 8'b00000000 ;
			15'h00004636 : data <= 8'b00000000 ;
			15'h00004637 : data <= 8'b00000000 ;
			15'h00004638 : data <= 8'b00000000 ;
			15'h00004639 : data <= 8'b00000000 ;
			15'h0000463A : data <= 8'b00000000 ;
			15'h0000463B : data <= 8'b00000000 ;
			15'h0000463C : data <= 8'b00000000 ;
			15'h0000463D : data <= 8'b00000000 ;
			15'h0000463E : data <= 8'b00000000 ;
			15'h0000463F : data <= 8'b00000000 ;
			15'h00004640 : data <= 8'b00000000 ;
			15'h00004641 : data <= 8'b00000000 ;
			15'h00004642 : data <= 8'b00000000 ;
			15'h00004643 : data <= 8'b00000000 ;
			15'h00004644 : data <= 8'b00000000 ;
			15'h00004645 : data <= 8'b00000000 ;
			15'h00004646 : data <= 8'b00000000 ;
			15'h00004647 : data <= 8'b00000000 ;
			15'h00004648 : data <= 8'b00000000 ;
			15'h00004649 : data <= 8'b00000000 ;
			15'h0000464A : data <= 8'b00000000 ;
			15'h0000464B : data <= 8'b00000000 ;
			15'h0000464C : data <= 8'b00000000 ;
			15'h0000464D : data <= 8'b00000000 ;
			15'h0000464E : data <= 8'b00000000 ;
			15'h0000464F : data <= 8'b00000000 ;
			15'h00004650 : data <= 8'b00000000 ;
			15'h00004651 : data <= 8'b00000000 ;
			15'h00004652 : data <= 8'b00000000 ;
			15'h00004653 : data <= 8'b00000000 ;
			15'h00004654 : data <= 8'b00000000 ;
			15'h00004655 : data <= 8'b00000000 ;
			15'h00004656 : data <= 8'b00000000 ;
			15'h00004657 : data <= 8'b00000000 ;
			15'h00004658 : data <= 8'b00000000 ;
			15'h00004659 : data <= 8'b00000000 ;
			15'h0000465A : data <= 8'b00000000 ;
			15'h0000465B : data <= 8'b00000000 ;
			15'h0000465C : data <= 8'b00000000 ;
			15'h0000465D : data <= 8'b00000000 ;
			15'h0000465E : data <= 8'b00000000 ;
			15'h0000465F : data <= 8'b00000000 ;
			15'h00004660 : data <= 8'b00000000 ;
			15'h00004661 : data <= 8'b00000000 ;
			15'h00004662 : data <= 8'b00000000 ;
			15'h00004663 : data <= 8'b00000000 ;
			15'h00004664 : data <= 8'b00000000 ;
			15'h00004665 : data <= 8'b00000000 ;
			15'h00004666 : data <= 8'b00000000 ;
			15'h00004667 : data <= 8'b00000000 ;
			15'h00004668 : data <= 8'b00000000 ;
			15'h00004669 : data <= 8'b00000000 ;
			15'h0000466A : data <= 8'b00000000 ;
			15'h0000466B : data <= 8'b00000000 ;
			15'h0000466C : data <= 8'b00000000 ;
			15'h0000466D : data <= 8'b00000000 ;
			15'h0000466E : data <= 8'b00000000 ;
			15'h0000466F : data <= 8'b00000000 ;
			15'h00004670 : data <= 8'b00000000 ;
			15'h00004671 : data <= 8'b00000000 ;
			15'h00004672 : data <= 8'b00000000 ;
			15'h00004673 : data <= 8'b00000000 ;
			15'h00004674 : data <= 8'b00000000 ;
			15'h00004675 : data <= 8'b00000000 ;
			15'h00004676 : data <= 8'b00000000 ;
			15'h00004677 : data <= 8'b00000000 ;
			15'h00004678 : data <= 8'b00000000 ;
			15'h00004679 : data <= 8'b00000000 ;
			15'h0000467A : data <= 8'b00000000 ;
			15'h0000467B : data <= 8'b00000000 ;
			15'h0000467C : data <= 8'b00000000 ;
			15'h0000467D : data <= 8'b00000000 ;
			15'h0000467E : data <= 8'b00000000 ;
			15'h0000467F : data <= 8'b00000000 ;
			15'h00004680 : data <= 8'b00000000 ;
			15'h00004681 : data <= 8'b00000000 ;
			15'h00004682 : data <= 8'b00000000 ;
			15'h00004683 : data <= 8'b00000000 ;
			15'h00004684 : data <= 8'b00000000 ;
			15'h00004685 : data <= 8'b00000000 ;
			15'h00004686 : data <= 8'b00000000 ;
			15'h00004687 : data <= 8'b00000000 ;
			15'h00004688 : data <= 8'b00000000 ;
			15'h00004689 : data <= 8'b00000000 ;
			15'h0000468A : data <= 8'b00000000 ;
			15'h0000468B : data <= 8'b00000000 ;
			15'h0000468C : data <= 8'b00000000 ;
			15'h0000468D : data <= 8'b00000000 ;
			15'h0000468E : data <= 8'b00000000 ;
			15'h0000468F : data <= 8'b00000000 ;
			15'h00004690 : data <= 8'b00000000 ;
			15'h00004691 : data <= 8'b00000000 ;
			15'h00004692 : data <= 8'b00000000 ;
			15'h00004693 : data <= 8'b00000000 ;
			15'h00004694 : data <= 8'b00000000 ;
			15'h00004695 : data <= 8'b00000000 ;
			15'h00004696 : data <= 8'b00000000 ;
			15'h00004697 : data <= 8'b00000000 ;
			15'h00004698 : data <= 8'b00000000 ;
			15'h00004699 : data <= 8'b00000000 ;
			15'h0000469A : data <= 8'b00000000 ;
			15'h0000469B : data <= 8'b00000000 ;
			15'h0000469C : data <= 8'b00000000 ;
			15'h0000469D : data <= 8'b00000000 ;
			15'h0000469E : data <= 8'b00000000 ;
			15'h0000469F : data <= 8'b00000000 ;
			15'h000046A0 : data <= 8'b00000000 ;
			15'h000046A1 : data <= 8'b00000000 ;
			15'h000046A2 : data <= 8'b00000000 ;
			15'h000046A3 : data <= 8'b00000000 ;
			15'h000046A4 : data <= 8'b00000000 ;
			15'h000046A5 : data <= 8'b00000000 ;
			15'h000046A6 : data <= 8'b00000000 ;
			15'h000046A7 : data <= 8'b00000000 ;
			15'h000046A8 : data <= 8'b00000000 ;
			15'h000046A9 : data <= 8'b00000000 ;
			15'h000046AA : data <= 8'b00000000 ;
			15'h000046AB : data <= 8'b00000000 ;
			15'h000046AC : data <= 8'b00000000 ;
			15'h000046AD : data <= 8'b00000000 ;
			15'h000046AE : data <= 8'b00000000 ;
			15'h000046AF : data <= 8'b00000000 ;
			15'h000046B0 : data <= 8'b00000000 ;
			15'h000046B1 : data <= 8'b00000000 ;
			15'h000046B2 : data <= 8'b00000000 ;
			15'h000046B3 : data <= 8'b00000000 ;
			15'h000046B4 : data <= 8'b00000000 ;
			15'h000046B5 : data <= 8'b00000000 ;
			15'h000046B6 : data <= 8'b00000000 ;
			15'h000046B7 : data <= 8'b00000000 ;
			15'h000046B8 : data <= 8'b00000000 ;
			15'h000046B9 : data <= 8'b00000000 ;
			15'h000046BA : data <= 8'b00000000 ;
			15'h000046BB : data <= 8'b00000000 ;
			15'h000046BC : data <= 8'b00000000 ;
			15'h000046BD : data <= 8'b00000000 ;
			15'h000046BE : data <= 8'b00000000 ;
			15'h000046BF : data <= 8'b00000000 ;
			15'h000046C0 : data <= 8'b00000000 ;
			15'h000046C1 : data <= 8'b00000000 ;
			15'h000046C2 : data <= 8'b00000000 ;
			15'h000046C3 : data <= 8'b00000000 ;
			15'h000046C4 : data <= 8'b00000000 ;
			15'h000046C5 : data <= 8'b00000000 ;
			15'h000046C6 : data <= 8'b00000000 ;
			15'h000046C7 : data <= 8'b00000000 ;
			15'h000046C8 : data <= 8'b00000000 ;
			15'h000046C9 : data <= 8'b00000000 ;
			15'h000046CA : data <= 8'b00000000 ;
			15'h000046CB : data <= 8'b00000000 ;
			15'h000046CC : data <= 8'b00000000 ;
			15'h000046CD : data <= 8'b00000000 ;
			15'h000046CE : data <= 8'b00000000 ;
			15'h000046CF : data <= 8'b00000000 ;
			15'h000046D0 : data <= 8'b00000000 ;
			15'h000046D1 : data <= 8'b00000000 ;
			15'h000046D2 : data <= 8'b00000000 ;
			15'h000046D3 : data <= 8'b00000000 ;
			15'h000046D4 : data <= 8'b00000000 ;
			15'h000046D5 : data <= 8'b00000000 ;
			15'h000046D6 : data <= 8'b00000000 ;
			15'h000046D7 : data <= 8'b00000000 ;
			15'h000046D8 : data <= 8'b00000000 ;
			15'h000046D9 : data <= 8'b00000000 ;
			15'h000046DA : data <= 8'b00000000 ;
			15'h000046DB : data <= 8'b00000000 ;
			15'h000046DC : data <= 8'b00000000 ;
			15'h000046DD : data <= 8'b00000000 ;
			15'h000046DE : data <= 8'b00000000 ;
			15'h000046DF : data <= 8'b00000000 ;
			15'h000046E0 : data <= 8'b00000000 ;
			15'h000046E1 : data <= 8'b00000000 ;
			15'h000046E2 : data <= 8'b00000000 ;
			15'h000046E3 : data <= 8'b00000000 ;
			15'h000046E4 : data <= 8'b00000000 ;
			15'h000046E5 : data <= 8'b00000000 ;
			15'h000046E6 : data <= 8'b00000000 ;
			15'h000046E7 : data <= 8'b00000000 ;
			15'h000046E8 : data <= 8'b00000000 ;
			15'h000046E9 : data <= 8'b00000000 ;
			15'h000046EA : data <= 8'b00000000 ;
			15'h000046EB : data <= 8'b00000000 ;
			15'h000046EC : data <= 8'b00000000 ;
			15'h000046ED : data <= 8'b00000000 ;
			15'h000046EE : data <= 8'b00000000 ;
			15'h000046EF : data <= 8'b00000000 ;
			15'h000046F0 : data <= 8'b00000000 ;
			15'h000046F1 : data <= 8'b00000000 ;
			15'h000046F2 : data <= 8'b00000000 ;
			15'h000046F3 : data <= 8'b00000000 ;
			15'h000046F4 : data <= 8'b00000000 ;
			15'h000046F5 : data <= 8'b00000000 ;
			15'h000046F6 : data <= 8'b00000000 ;
			15'h000046F7 : data <= 8'b00000000 ;
			15'h000046F8 : data <= 8'b00000000 ;
			15'h000046F9 : data <= 8'b00000000 ;
			15'h000046FA : data <= 8'b00000000 ;
			15'h000046FB : data <= 8'b00000000 ;
			15'h000046FC : data <= 8'b00000000 ;
			15'h000046FD : data <= 8'b00000000 ;
			15'h000046FE : data <= 8'b00000000 ;
			15'h000046FF : data <= 8'b00000000 ;
			15'h00004700 : data <= 8'b00000000 ;
			15'h00004701 : data <= 8'b00000000 ;
			15'h00004702 : data <= 8'b00000000 ;
			15'h00004703 : data <= 8'b00000000 ;
			15'h00004704 : data <= 8'b00000000 ;
			15'h00004705 : data <= 8'b00000000 ;
			15'h00004706 : data <= 8'b00000000 ;
			15'h00004707 : data <= 8'b00000000 ;
			15'h00004708 : data <= 8'b00000000 ;
			15'h00004709 : data <= 8'b00000000 ;
			15'h0000470A : data <= 8'b00000000 ;
			15'h0000470B : data <= 8'b00000000 ;
			15'h0000470C : data <= 8'b00000000 ;
			15'h0000470D : data <= 8'b00000000 ;
			15'h0000470E : data <= 8'b00000000 ;
			15'h0000470F : data <= 8'b00000000 ;
			15'h00004710 : data <= 8'b00000000 ;
			15'h00004711 : data <= 8'b00000000 ;
			15'h00004712 : data <= 8'b00000000 ;
			15'h00004713 : data <= 8'b00000000 ;
			15'h00004714 : data <= 8'b00000000 ;
			15'h00004715 : data <= 8'b00000000 ;
			15'h00004716 : data <= 8'b00000000 ;
			15'h00004717 : data <= 8'b00000000 ;
			15'h00004718 : data <= 8'b00000000 ;
			15'h00004719 : data <= 8'b00000000 ;
			15'h0000471A : data <= 8'b00000000 ;
			15'h0000471B : data <= 8'b00000000 ;
			15'h0000471C : data <= 8'b00000000 ;
			15'h0000471D : data <= 8'b00000000 ;
			15'h0000471E : data <= 8'b00000000 ;
			15'h0000471F : data <= 8'b00000000 ;
			15'h00004720 : data <= 8'b00000000 ;
			15'h00004721 : data <= 8'b00000000 ;
			15'h00004722 : data <= 8'b00000000 ;
			15'h00004723 : data <= 8'b00000000 ;
			15'h00004724 : data <= 8'b00000000 ;
			15'h00004725 : data <= 8'b00000000 ;
			15'h00004726 : data <= 8'b00000000 ;
			15'h00004727 : data <= 8'b00000000 ;
			15'h00004728 : data <= 8'b00000000 ;
			15'h00004729 : data <= 8'b00000000 ;
			15'h0000472A : data <= 8'b00000000 ;
			15'h0000472B : data <= 8'b00000000 ;
			15'h0000472C : data <= 8'b00000000 ;
			15'h0000472D : data <= 8'b00000000 ;
			15'h0000472E : data <= 8'b00000000 ;
			15'h0000472F : data <= 8'b00000000 ;
			15'h00004730 : data <= 8'b00000000 ;
			15'h00004731 : data <= 8'b00000000 ;
			15'h00004732 : data <= 8'b00000000 ;
			15'h00004733 : data <= 8'b00000000 ;
			15'h00004734 : data <= 8'b00000000 ;
			15'h00004735 : data <= 8'b00000000 ;
			15'h00004736 : data <= 8'b00000000 ;
			15'h00004737 : data <= 8'b00000000 ;
			15'h00004738 : data <= 8'b00000000 ;
			15'h00004739 : data <= 8'b00000000 ;
			15'h0000473A : data <= 8'b00000000 ;
			15'h0000473B : data <= 8'b00000000 ;
			15'h0000473C : data <= 8'b00000000 ;
			15'h0000473D : data <= 8'b00000000 ;
			15'h0000473E : data <= 8'b00000000 ;
			15'h0000473F : data <= 8'b00000000 ;
			15'h00004740 : data <= 8'b00000000 ;
			15'h00004741 : data <= 8'b00000000 ;
			15'h00004742 : data <= 8'b00000000 ;
			15'h00004743 : data <= 8'b00000000 ;
			15'h00004744 : data <= 8'b00000000 ;
			15'h00004745 : data <= 8'b00000000 ;
			15'h00004746 : data <= 8'b00000000 ;
			15'h00004747 : data <= 8'b00000000 ;
			15'h00004748 : data <= 8'b00000000 ;
			15'h00004749 : data <= 8'b00000000 ;
			15'h0000474A : data <= 8'b00000000 ;
			15'h0000474B : data <= 8'b00000000 ;
			15'h0000474C : data <= 8'b00000000 ;
			15'h0000474D : data <= 8'b00000000 ;
			15'h0000474E : data <= 8'b00000000 ;
			15'h0000474F : data <= 8'b00000000 ;
			15'h00004750 : data <= 8'b00000000 ;
			15'h00004751 : data <= 8'b00000000 ;
			15'h00004752 : data <= 8'b00000000 ;
			15'h00004753 : data <= 8'b00000000 ;
			15'h00004754 : data <= 8'b00000000 ;
			15'h00004755 : data <= 8'b00000000 ;
			15'h00004756 : data <= 8'b00000000 ;
			15'h00004757 : data <= 8'b00000000 ;
			15'h00004758 : data <= 8'b00000000 ;
			15'h00004759 : data <= 8'b00000000 ;
			15'h0000475A : data <= 8'b00000000 ;
			15'h0000475B : data <= 8'b00000000 ;
			15'h0000475C : data <= 8'b00000000 ;
			15'h0000475D : data <= 8'b00000000 ;
			15'h0000475E : data <= 8'b00000000 ;
			15'h0000475F : data <= 8'b00000000 ;
			15'h00004760 : data <= 8'b00000000 ;
			15'h00004761 : data <= 8'b00000000 ;
			15'h00004762 : data <= 8'b00000000 ;
			15'h00004763 : data <= 8'b00000000 ;
			15'h00004764 : data <= 8'b00000000 ;
			15'h00004765 : data <= 8'b00000000 ;
			15'h00004766 : data <= 8'b00000000 ;
			15'h00004767 : data <= 8'b00000000 ;
			15'h00004768 : data <= 8'b00000000 ;
			15'h00004769 : data <= 8'b00000000 ;
			15'h0000476A : data <= 8'b00000000 ;
			15'h0000476B : data <= 8'b00000000 ;
			15'h0000476C : data <= 8'b00000000 ;
			15'h0000476D : data <= 8'b00000000 ;
			15'h0000476E : data <= 8'b00000000 ;
			15'h0000476F : data <= 8'b00000000 ;
			15'h00004770 : data <= 8'b00000000 ;
			15'h00004771 : data <= 8'b00000000 ;
			15'h00004772 : data <= 8'b00000000 ;
			15'h00004773 : data <= 8'b00000000 ;
			15'h00004774 : data <= 8'b00000000 ;
			15'h00004775 : data <= 8'b00000000 ;
			15'h00004776 : data <= 8'b00000000 ;
			15'h00004777 : data <= 8'b00000000 ;
			15'h00004778 : data <= 8'b00000000 ;
			15'h00004779 : data <= 8'b00000000 ;
			15'h0000477A : data <= 8'b00000000 ;
			15'h0000477B : data <= 8'b00000000 ;
			15'h0000477C : data <= 8'b00000000 ;
			15'h0000477D : data <= 8'b00000000 ;
			15'h0000477E : data <= 8'b00000000 ;
			15'h0000477F : data <= 8'b00000000 ;
			15'h00004780 : data <= 8'b00000000 ;
			15'h00004781 : data <= 8'b00000000 ;
			15'h00004782 : data <= 8'b00000000 ;
			15'h00004783 : data <= 8'b00000000 ;
			15'h00004784 : data <= 8'b00000000 ;
			15'h00004785 : data <= 8'b00000000 ;
			15'h00004786 : data <= 8'b00000000 ;
			15'h00004787 : data <= 8'b00000000 ;
			15'h00004788 : data <= 8'b00000000 ;
			15'h00004789 : data <= 8'b00000000 ;
			15'h0000478A : data <= 8'b00000000 ;
			15'h0000478B : data <= 8'b00000000 ;
			15'h0000478C : data <= 8'b00000000 ;
			15'h0000478D : data <= 8'b00000000 ;
			15'h0000478E : data <= 8'b00000000 ;
			15'h0000478F : data <= 8'b00000000 ;
			15'h00004790 : data <= 8'b00000000 ;
			15'h00004791 : data <= 8'b00000000 ;
			15'h00004792 : data <= 8'b00000000 ;
			15'h00004793 : data <= 8'b00000000 ;
			15'h00004794 : data <= 8'b00000000 ;
			15'h00004795 : data <= 8'b00000000 ;
			15'h00004796 : data <= 8'b00000000 ;
			15'h00004797 : data <= 8'b00000000 ;
			15'h00004798 : data <= 8'b00000000 ;
			15'h00004799 : data <= 8'b00000000 ;
			15'h0000479A : data <= 8'b00000000 ;
			15'h0000479B : data <= 8'b00000000 ;
			15'h0000479C : data <= 8'b00000000 ;
			15'h0000479D : data <= 8'b00000000 ;
			15'h0000479E : data <= 8'b00000000 ;
			15'h0000479F : data <= 8'b00000000 ;
			15'h000047A0 : data <= 8'b00000000 ;
			15'h000047A1 : data <= 8'b00000000 ;
			15'h000047A2 : data <= 8'b00000000 ;
			15'h000047A3 : data <= 8'b00000000 ;
			15'h000047A4 : data <= 8'b00000000 ;
			15'h000047A5 : data <= 8'b00000000 ;
			15'h000047A6 : data <= 8'b00000000 ;
			15'h000047A7 : data <= 8'b00000000 ;
			15'h000047A8 : data <= 8'b00000000 ;
			15'h000047A9 : data <= 8'b00000000 ;
			15'h000047AA : data <= 8'b00000000 ;
			15'h000047AB : data <= 8'b00000000 ;
			15'h000047AC : data <= 8'b00000000 ;
			15'h000047AD : data <= 8'b00000000 ;
			15'h000047AE : data <= 8'b00000000 ;
			15'h000047AF : data <= 8'b00000000 ;
			15'h000047B0 : data <= 8'b00000000 ;
			15'h000047B1 : data <= 8'b00000000 ;
			15'h000047B2 : data <= 8'b00000000 ;
			15'h000047B3 : data <= 8'b00000000 ;
			15'h000047B4 : data <= 8'b00000000 ;
			15'h000047B5 : data <= 8'b00000000 ;
			15'h000047B6 : data <= 8'b00000000 ;
			15'h000047B7 : data <= 8'b00000000 ;
			15'h000047B8 : data <= 8'b00000000 ;
			15'h000047B9 : data <= 8'b00000000 ;
			15'h000047BA : data <= 8'b00000000 ;
			15'h000047BB : data <= 8'b00000000 ;
			15'h000047BC : data <= 8'b00000000 ;
			15'h000047BD : data <= 8'b00000000 ;
			15'h000047BE : data <= 8'b00000000 ;
			15'h000047BF : data <= 8'b00000000 ;
			15'h000047C0 : data <= 8'b00000000 ;
			15'h000047C1 : data <= 8'b00000000 ;
			15'h000047C2 : data <= 8'b00000000 ;
			15'h000047C3 : data <= 8'b00000000 ;
			15'h000047C4 : data <= 8'b00000000 ;
			15'h000047C5 : data <= 8'b00000000 ;
			15'h000047C6 : data <= 8'b00000000 ;
			15'h000047C7 : data <= 8'b00000000 ;
			15'h000047C8 : data <= 8'b00000000 ;
			15'h000047C9 : data <= 8'b00000000 ;
			15'h000047CA : data <= 8'b00000000 ;
			15'h000047CB : data <= 8'b00000000 ;
			15'h000047CC : data <= 8'b00000000 ;
			15'h000047CD : data <= 8'b00000000 ;
			15'h000047CE : data <= 8'b00000000 ;
			15'h000047CF : data <= 8'b00000000 ;
			15'h000047D0 : data <= 8'b00000000 ;
			15'h000047D1 : data <= 8'b00000000 ;
			15'h000047D2 : data <= 8'b00000000 ;
			15'h000047D3 : data <= 8'b00000000 ;
			15'h000047D4 : data <= 8'b00000000 ;
			15'h000047D5 : data <= 8'b00000000 ;
			15'h000047D6 : data <= 8'b00000000 ;
			15'h000047D7 : data <= 8'b00000000 ;
			15'h000047D8 : data <= 8'b00000000 ;
			15'h000047D9 : data <= 8'b00000000 ;
			15'h000047DA : data <= 8'b00000000 ;
			15'h000047DB : data <= 8'b00000000 ;
			15'h000047DC : data <= 8'b00000000 ;
			15'h000047DD : data <= 8'b00000000 ;
			15'h000047DE : data <= 8'b00000000 ;
			15'h000047DF : data <= 8'b00000000 ;
			15'h000047E0 : data <= 8'b00000000 ;
			15'h000047E1 : data <= 8'b00000000 ;
			15'h000047E2 : data <= 8'b00000000 ;
			15'h000047E3 : data <= 8'b00000000 ;
			15'h000047E4 : data <= 8'b00000000 ;
			15'h000047E5 : data <= 8'b00000000 ;
			15'h000047E6 : data <= 8'b00000000 ;
			15'h000047E7 : data <= 8'b00000000 ;
			15'h000047E8 : data <= 8'b00000000 ;
			15'h000047E9 : data <= 8'b00000000 ;
			15'h000047EA : data <= 8'b00000000 ;
			15'h000047EB : data <= 8'b00000000 ;
			15'h000047EC : data <= 8'b00000000 ;
			15'h000047ED : data <= 8'b00000000 ;
			15'h000047EE : data <= 8'b00000000 ;
			15'h000047EF : data <= 8'b00000000 ;
			15'h000047F0 : data <= 8'b00000000 ;
			15'h000047F1 : data <= 8'b00000000 ;
			15'h000047F2 : data <= 8'b00000000 ;
			15'h000047F3 : data <= 8'b00000000 ;
			15'h000047F4 : data <= 8'b00000000 ;
			15'h000047F5 : data <= 8'b00000000 ;
			15'h000047F6 : data <= 8'b00000000 ;
			15'h000047F7 : data <= 8'b00000000 ;
			15'h000047F8 : data <= 8'b00000000 ;
			15'h000047F9 : data <= 8'b00000000 ;
			15'h000047FA : data <= 8'b00000000 ;
			15'h000047FB : data <= 8'b00000000 ;
			15'h000047FC : data <= 8'b00000000 ;
			15'h000047FD : data <= 8'b00000000 ;
			15'h000047FE : data <= 8'b00000000 ;
			15'h000047FF : data <= 8'b00000000 ;
			15'h00004800 : data <= 8'b00000000 ;
			15'h00004801 : data <= 8'b00000000 ;
			15'h00004802 : data <= 8'b00000000 ;
			15'h00004803 : data <= 8'b00000000 ;
			15'h00004804 : data <= 8'b00000000 ;
			15'h00004805 : data <= 8'b00000000 ;
			15'h00004806 : data <= 8'b00000000 ;
			15'h00004807 : data <= 8'b00000000 ;
			15'h00004808 : data <= 8'b00000000 ;
			15'h00004809 : data <= 8'b00000000 ;
			15'h0000480A : data <= 8'b00000000 ;
			15'h0000480B : data <= 8'b00000000 ;
			15'h0000480C : data <= 8'b00000000 ;
			15'h0000480D : data <= 8'b00000000 ;
			15'h0000480E : data <= 8'b00000000 ;
			15'h0000480F : data <= 8'b00000000 ;
			15'h00004810 : data <= 8'b00000000 ;
			15'h00004811 : data <= 8'b00000000 ;
			15'h00004812 : data <= 8'b00000000 ;
			15'h00004813 : data <= 8'b00000000 ;
			15'h00004814 : data <= 8'b00000000 ;
			15'h00004815 : data <= 8'b00000000 ;
			15'h00004816 : data <= 8'b00000000 ;
			15'h00004817 : data <= 8'b00000000 ;
			15'h00004818 : data <= 8'b00000000 ;
			15'h00004819 : data <= 8'b00000000 ;
			15'h0000481A : data <= 8'b00000000 ;
			15'h0000481B : data <= 8'b00000000 ;
			15'h0000481C : data <= 8'b00000000 ;
			15'h0000481D : data <= 8'b00000000 ;
			15'h0000481E : data <= 8'b00000000 ;
			15'h0000481F : data <= 8'b00000000 ;
			15'h00004820 : data <= 8'b00000000 ;
			15'h00004821 : data <= 8'b00000000 ;
			15'h00004822 : data <= 8'b00000000 ;
			15'h00004823 : data <= 8'b00000000 ;
			15'h00004824 : data <= 8'b00000000 ;
			15'h00004825 : data <= 8'b00000000 ;
			15'h00004826 : data <= 8'b00000000 ;
			15'h00004827 : data <= 8'b00000000 ;
			15'h00004828 : data <= 8'b00000000 ;
			15'h00004829 : data <= 8'b00000000 ;
			15'h0000482A : data <= 8'b00000000 ;
			15'h0000482B : data <= 8'b00000000 ;
			15'h0000482C : data <= 8'b00000000 ;
			15'h0000482D : data <= 8'b00000000 ;
			15'h0000482E : data <= 8'b00000000 ;
			15'h0000482F : data <= 8'b00000000 ;
			15'h00004830 : data <= 8'b00000000 ;
			15'h00004831 : data <= 8'b00000000 ;
			15'h00004832 : data <= 8'b00000000 ;
			15'h00004833 : data <= 8'b00000000 ;
			15'h00004834 : data <= 8'b00000000 ;
			15'h00004835 : data <= 8'b00000000 ;
			15'h00004836 : data <= 8'b00000000 ;
			15'h00004837 : data <= 8'b00000000 ;
			15'h00004838 : data <= 8'b00000000 ;
			15'h00004839 : data <= 8'b00000000 ;
			15'h0000483A : data <= 8'b00000000 ;
			15'h0000483B : data <= 8'b00000000 ;
			15'h0000483C : data <= 8'b00000000 ;
			15'h0000483D : data <= 8'b00000000 ;
			15'h0000483E : data <= 8'b00000000 ;
			15'h0000483F : data <= 8'b00000000 ;
			15'h00004840 : data <= 8'b00000000 ;
			15'h00004841 : data <= 8'b00000000 ;
			15'h00004842 : data <= 8'b00000000 ;
			15'h00004843 : data <= 8'b00000000 ;
			15'h00004844 : data <= 8'b00000000 ;
			15'h00004845 : data <= 8'b00000000 ;
			15'h00004846 : data <= 8'b00000000 ;
			15'h00004847 : data <= 8'b00000000 ;
			15'h00004848 : data <= 8'b00000000 ;
			15'h00004849 : data <= 8'b00000000 ;
			15'h0000484A : data <= 8'b00000000 ;
			15'h0000484B : data <= 8'b00000000 ;
			15'h0000484C : data <= 8'b00000000 ;
			15'h0000484D : data <= 8'b00000000 ;
			15'h0000484E : data <= 8'b00000000 ;
			15'h0000484F : data <= 8'b00000000 ;
			15'h00004850 : data <= 8'b00000000 ;
			15'h00004851 : data <= 8'b00000000 ;
			15'h00004852 : data <= 8'b00000000 ;
			15'h00004853 : data <= 8'b00000000 ;
			15'h00004854 : data <= 8'b00000000 ;
			15'h00004855 : data <= 8'b00000000 ;
			15'h00004856 : data <= 8'b00000000 ;
			15'h00004857 : data <= 8'b00000000 ;
			15'h00004858 : data <= 8'b00000000 ;
			15'h00004859 : data <= 8'b00000000 ;
			15'h0000485A : data <= 8'b00000000 ;
			15'h0000485B : data <= 8'b00000000 ;
			15'h0000485C : data <= 8'b00000000 ;
			15'h0000485D : data <= 8'b00000000 ;
			15'h0000485E : data <= 8'b00000000 ;
			15'h0000485F : data <= 8'b00000000 ;
			15'h00004860 : data <= 8'b00000000 ;
			15'h00004861 : data <= 8'b00000000 ;
			15'h00004862 : data <= 8'b00000000 ;
			15'h00004863 : data <= 8'b00000000 ;
			15'h00004864 : data <= 8'b00000000 ;
			15'h00004865 : data <= 8'b00000000 ;
			15'h00004866 : data <= 8'b00000000 ;
			15'h00004867 : data <= 8'b00000000 ;
			15'h00004868 : data <= 8'b00000000 ;
			15'h00004869 : data <= 8'b00000000 ;
			15'h0000486A : data <= 8'b00000000 ;
			15'h0000486B : data <= 8'b00000000 ;
			15'h0000486C : data <= 8'b00000000 ;
			15'h0000486D : data <= 8'b00000000 ;
			15'h0000486E : data <= 8'b00000000 ;
			15'h0000486F : data <= 8'b00000000 ;
			15'h00004870 : data <= 8'b00000000 ;
			15'h00004871 : data <= 8'b00000000 ;
			15'h00004872 : data <= 8'b00000000 ;
			15'h00004873 : data <= 8'b00000000 ;
			15'h00004874 : data <= 8'b00000000 ;
			15'h00004875 : data <= 8'b00000000 ;
			15'h00004876 : data <= 8'b00000000 ;
			15'h00004877 : data <= 8'b00000000 ;
			15'h00004878 : data <= 8'b00000000 ;
			15'h00004879 : data <= 8'b00000000 ;
			15'h0000487A : data <= 8'b00000000 ;
			15'h0000487B : data <= 8'b00000000 ;
			15'h0000487C : data <= 8'b00000000 ;
			15'h0000487D : data <= 8'b00000000 ;
			15'h0000487E : data <= 8'b00000000 ;
			15'h0000487F : data <= 8'b00000000 ;
			15'h00004880 : data <= 8'b00000000 ;
			15'h00004881 : data <= 8'b00000000 ;
			15'h00004882 : data <= 8'b00000000 ;
			15'h00004883 : data <= 8'b00000000 ;
			15'h00004884 : data <= 8'b00000000 ;
			15'h00004885 : data <= 8'b00000000 ;
			15'h00004886 : data <= 8'b00000000 ;
			15'h00004887 : data <= 8'b00000000 ;
			15'h00004888 : data <= 8'b00000000 ;
			15'h00004889 : data <= 8'b00000000 ;
			15'h0000488A : data <= 8'b00000000 ;
			15'h0000488B : data <= 8'b00000000 ;
			15'h0000488C : data <= 8'b00000000 ;
			15'h0000488D : data <= 8'b00000000 ;
			15'h0000488E : data <= 8'b00000000 ;
			15'h0000488F : data <= 8'b00000000 ;
			15'h00004890 : data <= 8'b00000000 ;
			15'h00004891 : data <= 8'b00000000 ;
			15'h00004892 : data <= 8'b00000000 ;
			15'h00004893 : data <= 8'b00000000 ;
			15'h00004894 : data <= 8'b00000000 ;
			15'h00004895 : data <= 8'b00000000 ;
			15'h00004896 : data <= 8'b00000000 ;
			15'h00004897 : data <= 8'b00000000 ;
			15'h00004898 : data <= 8'b00000000 ;
			15'h00004899 : data <= 8'b00000000 ;
			15'h0000489A : data <= 8'b00000000 ;
			15'h0000489B : data <= 8'b00000000 ;
			15'h0000489C : data <= 8'b00000000 ;
			15'h0000489D : data <= 8'b00000000 ;
			15'h0000489E : data <= 8'b00000000 ;
			15'h0000489F : data <= 8'b00000000 ;
			15'h000048A0 : data <= 8'b00000000 ;
			15'h000048A1 : data <= 8'b00000000 ;
			15'h000048A2 : data <= 8'b00000000 ;
			15'h000048A3 : data <= 8'b00000000 ;
			15'h000048A4 : data <= 8'b00000000 ;
			15'h000048A5 : data <= 8'b00000000 ;
			15'h000048A6 : data <= 8'b00000000 ;
			15'h000048A7 : data <= 8'b00000000 ;
			15'h000048A8 : data <= 8'b00000000 ;
			15'h000048A9 : data <= 8'b00000000 ;
			15'h000048AA : data <= 8'b00000000 ;
			15'h000048AB : data <= 8'b00000000 ;
			15'h000048AC : data <= 8'b00000000 ;
			15'h000048AD : data <= 8'b00000000 ;
			15'h000048AE : data <= 8'b00000000 ;
			15'h000048AF : data <= 8'b00000000 ;
			15'h000048B0 : data <= 8'b00000000 ;
			15'h000048B1 : data <= 8'b00000000 ;
			15'h000048B2 : data <= 8'b00000000 ;
			15'h000048B3 : data <= 8'b00000000 ;
			15'h000048B4 : data <= 8'b00000000 ;
			15'h000048B5 : data <= 8'b00000000 ;
			15'h000048B6 : data <= 8'b00000000 ;
			15'h000048B7 : data <= 8'b00000000 ;
			15'h000048B8 : data <= 8'b00000000 ;
			15'h000048B9 : data <= 8'b00000000 ;
			15'h000048BA : data <= 8'b00000000 ;
			15'h000048BB : data <= 8'b00000000 ;
			15'h000048BC : data <= 8'b00000000 ;
			15'h000048BD : data <= 8'b00000000 ;
			15'h000048BE : data <= 8'b00000000 ;
			15'h000048BF : data <= 8'b00000000 ;
			15'h000048C0 : data <= 8'b00000000 ;
			15'h000048C1 : data <= 8'b00000000 ;
			15'h000048C2 : data <= 8'b00000000 ;
			15'h000048C3 : data <= 8'b00000000 ;
			15'h000048C4 : data <= 8'b00000000 ;
			15'h000048C5 : data <= 8'b00000000 ;
			15'h000048C6 : data <= 8'b00000000 ;
			15'h000048C7 : data <= 8'b00000000 ;
			15'h000048C8 : data <= 8'b00000000 ;
			15'h000048C9 : data <= 8'b00000000 ;
			15'h000048CA : data <= 8'b00000000 ;
			15'h000048CB : data <= 8'b00000000 ;
			15'h000048CC : data <= 8'b00000000 ;
			15'h000048CD : data <= 8'b00000000 ;
			15'h000048CE : data <= 8'b00000000 ;
			15'h000048CF : data <= 8'b00000000 ;
			15'h000048D0 : data <= 8'b00000000 ;
			15'h000048D1 : data <= 8'b00000000 ;
			15'h000048D2 : data <= 8'b00000000 ;
			15'h000048D3 : data <= 8'b00000000 ;
			15'h000048D4 : data <= 8'b00000000 ;
			15'h000048D5 : data <= 8'b00000000 ;
			15'h000048D6 : data <= 8'b00000000 ;
			15'h000048D7 : data <= 8'b00000000 ;
			15'h000048D8 : data <= 8'b00000000 ;
			15'h000048D9 : data <= 8'b00000000 ;
			15'h000048DA : data <= 8'b00000000 ;
			15'h000048DB : data <= 8'b00000000 ;
			15'h000048DC : data <= 8'b00000000 ;
			15'h000048DD : data <= 8'b00000000 ;
			15'h000048DE : data <= 8'b00000000 ;
			15'h000048DF : data <= 8'b00000000 ;
			15'h000048E0 : data <= 8'b00000000 ;
			15'h000048E1 : data <= 8'b00000000 ;
			15'h000048E2 : data <= 8'b00000000 ;
			15'h000048E3 : data <= 8'b00000000 ;
			15'h000048E4 : data <= 8'b00000000 ;
			15'h000048E5 : data <= 8'b00000000 ;
			15'h000048E6 : data <= 8'b00000000 ;
			15'h000048E7 : data <= 8'b00000000 ;
			15'h000048E8 : data <= 8'b00000000 ;
			15'h000048E9 : data <= 8'b00000000 ;
			15'h000048EA : data <= 8'b00000000 ;
			15'h000048EB : data <= 8'b00000000 ;
			15'h000048EC : data <= 8'b00000000 ;
			15'h000048ED : data <= 8'b00000000 ;
			15'h000048EE : data <= 8'b00000000 ;
			15'h000048EF : data <= 8'b00000000 ;
			15'h000048F0 : data <= 8'b00000000 ;
			15'h000048F1 : data <= 8'b00000000 ;
			15'h000048F2 : data <= 8'b00000000 ;
			15'h000048F3 : data <= 8'b00000000 ;
			15'h000048F4 : data <= 8'b00000000 ;
			15'h000048F5 : data <= 8'b00000000 ;
			15'h000048F6 : data <= 8'b00000000 ;
			15'h000048F7 : data <= 8'b00000000 ;
			15'h000048F8 : data <= 8'b00000000 ;
			15'h000048F9 : data <= 8'b00000000 ;
			15'h000048FA : data <= 8'b00000000 ;
			15'h000048FB : data <= 8'b00000000 ;
			15'h000048FC : data <= 8'b00000000 ;
			15'h000048FD : data <= 8'b00000000 ;
			15'h000048FE : data <= 8'b00000000 ;
			15'h000048FF : data <= 8'b00000000 ;
			15'h00004900 : data <= 8'b00000000 ;
			15'h00004901 : data <= 8'b00000000 ;
			15'h00004902 : data <= 8'b00000000 ;
			15'h00004903 : data <= 8'b00000000 ;
			15'h00004904 : data <= 8'b00000000 ;
			15'h00004905 : data <= 8'b00000000 ;
			15'h00004906 : data <= 8'b00000000 ;
			15'h00004907 : data <= 8'b00000000 ;
			15'h00004908 : data <= 8'b00000000 ;
			15'h00004909 : data <= 8'b00000000 ;
			15'h0000490A : data <= 8'b00000000 ;
			15'h0000490B : data <= 8'b00000000 ;
			15'h0000490C : data <= 8'b00000000 ;
			15'h0000490D : data <= 8'b00000000 ;
			15'h0000490E : data <= 8'b00000000 ;
			15'h0000490F : data <= 8'b00000000 ;
			15'h00004910 : data <= 8'b00000000 ;
			15'h00004911 : data <= 8'b00000000 ;
			15'h00004912 : data <= 8'b00000000 ;
			15'h00004913 : data <= 8'b00000000 ;
			15'h00004914 : data <= 8'b00000000 ;
			15'h00004915 : data <= 8'b00000000 ;
			15'h00004916 : data <= 8'b00000000 ;
			15'h00004917 : data <= 8'b00000000 ;
			15'h00004918 : data <= 8'b00000000 ;
			15'h00004919 : data <= 8'b00000000 ;
			15'h0000491A : data <= 8'b00000000 ;
			15'h0000491B : data <= 8'b00000000 ;
			15'h0000491C : data <= 8'b00000000 ;
			15'h0000491D : data <= 8'b00000000 ;
			15'h0000491E : data <= 8'b00000000 ;
			15'h0000491F : data <= 8'b00000000 ;
			15'h00004920 : data <= 8'b00000000 ;
			15'h00004921 : data <= 8'b00000000 ;
			15'h00004922 : data <= 8'b00000000 ;
			15'h00004923 : data <= 8'b00000000 ;
			15'h00004924 : data <= 8'b00000000 ;
			15'h00004925 : data <= 8'b00000000 ;
			15'h00004926 : data <= 8'b00000000 ;
			15'h00004927 : data <= 8'b00000000 ;
			15'h00004928 : data <= 8'b00000000 ;
			15'h00004929 : data <= 8'b00000000 ;
			15'h0000492A : data <= 8'b00000000 ;
			15'h0000492B : data <= 8'b00000000 ;
			15'h0000492C : data <= 8'b00000000 ;
			15'h0000492D : data <= 8'b00000000 ;
			15'h0000492E : data <= 8'b00000000 ;
			15'h0000492F : data <= 8'b00000000 ;
			15'h00004930 : data <= 8'b00000000 ;
			15'h00004931 : data <= 8'b00000000 ;
			15'h00004932 : data <= 8'b00000000 ;
			15'h00004933 : data <= 8'b00000000 ;
			15'h00004934 : data <= 8'b00000000 ;
			15'h00004935 : data <= 8'b00000000 ;
			15'h00004936 : data <= 8'b00000000 ;
			15'h00004937 : data <= 8'b00000000 ;
			15'h00004938 : data <= 8'b00000000 ;
			15'h00004939 : data <= 8'b00000000 ;
			15'h0000493A : data <= 8'b00000000 ;
			15'h0000493B : data <= 8'b00000000 ;
			15'h0000493C : data <= 8'b00000000 ;
			15'h0000493D : data <= 8'b00000000 ;
			15'h0000493E : data <= 8'b00000000 ;
			15'h0000493F : data <= 8'b00000000 ;
			15'h00004940 : data <= 8'b00000000 ;
			15'h00004941 : data <= 8'b00000000 ;
			15'h00004942 : data <= 8'b00000000 ;
			15'h00004943 : data <= 8'b00000000 ;
			15'h00004944 : data <= 8'b00000000 ;
			15'h00004945 : data <= 8'b00000000 ;
			15'h00004946 : data <= 8'b00000000 ;
			15'h00004947 : data <= 8'b00000000 ;
			15'h00004948 : data <= 8'b00000000 ;
			15'h00004949 : data <= 8'b00000000 ;
			15'h0000494A : data <= 8'b00000000 ;
			15'h0000494B : data <= 8'b00000000 ;
			15'h0000494C : data <= 8'b00000000 ;
			15'h0000494D : data <= 8'b00000000 ;
			15'h0000494E : data <= 8'b00000000 ;
			15'h0000494F : data <= 8'b00000000 ;
			15'h00004950 : data <= 8'b00000000 ;
			15'h00004951 : data <= 8'b00000000 ;
			15'h00004952 : data <= 8'b00000000 ;
			15'h00004953 : data <= 8'b00000000 ;
			15'h00004954 : data <= 8'b00000000 ;
			15'h00004955 : data <= 8'b00000000 ;
			15'h00004956 : data <= 8'b00000000 ;
			15'h00004957 : data <= 8'b00000000 ;
			15'h00004958 : data <= 8'b00000000 ;
			15'h00004959 : data <= 8'b00000000 ;
			15'h0000495A : data <= 8'b00000000 ;
			15'h0000495B : data <= 8'b00000000 ;
			15'h0000495C : data <= 8'b00000000 ;
			15'h0000495D : data <= 8'b00000000 ;
			15'h0000495E : data <= 8'b00000000 ;
			15'h0000495F : data <= 8'b00000000 ;
			15'h00004960 : data <= 8'b00000000 ;
			15'h00004961 : data <= 8'b00000000 ;
			15'h00004962 : data <= 8'b00000000 ;
			15'h00004963 : data <= 8'b00000000 ;
			15'h00004964 : data <= 8'b00000000 ;
			15'h00004965 : data <= 8'b00000000 ;
			15'h00004966 : data <= 8'b00000000 ;
			15'h00004967 : data <= 8'b00000000 ;
			15'h00004968 : data <= 8'b00000000 ;
			15'h00004969 : data <= 8'b00000000 ;
			15'h0000496A : data <= 8'b00000000 ;
			15'h0000496B : data <= 8'b00000000 ;
			15'h0000496C : data <= 8'b00000000 ;
			15'h0000496D : data <= 8'b00000000 ;
			15'h0000496E : data <= 8'b00000000 ;
			15'h0000496F : data <= 8'b00000000 ;
			15'h00004970 : data <= 8'b00000000 ;
			15'h00004971 : data <= 8'b00000000 ;
			15'h00004972 : data <= 8'b00000000 ;
			15'h00004973 : data <= 8'b00000000 ;
			15'h00004974 : data <= 8'b00000000 ;
			15'h00004975 : data <= 8'b00000000 ;
			15'h00004976 : data <= 8'b00000000 ;
			15'h00004977 : data <= 8'b00000000 ;
			15'h00004978 : data <= 8'b00000000 ;
			15'h00004979 : data <= 8'b00000000 ;
			15'h0000497A : data <= 8'b00000000 ;
			15'h0000497B : data <= 8'b00000000 ;
			15'h0000497C : data <= 8'b00000000 ;
			15'h0000497D : data <= 8'b00000000 ;
			15'h0000497E : data <= 8'b00000000 ;
			15'h0000497F : data <= 8'b00000000 ;
			15'h00004980 : data <= 8'b00000000 ;
			15'h00004981 : data <= 8'b00000000 ;
			15'h00004982 : data <= 8'b00000000 ;
			15'h00004983 : data <= 8'b00000000 ;
			15'h00004984 : data <= 8'b00000000 ;
			15'h00004985 : data <= 8'b00000000 ;
			15'h00004986 : data <= 8'b00000000 ;
			15'h00004987 : data <= 8'b00000000 ;
			15'h00004988 : data <= 8'b00000000 ;
			15'h00004989 : data <= 8'b00000000 ;
			15'h0000498A : data <= 8'b00000000 ;
			15'h0000498B : data <= 8'b00000000 ;
			15'h0000498C : data <= 8'b00000000 ;
			15'h0000498D : data <= 8'b00000000 ;
			15'h0000498E : data <= 8'b00000000 ;
			15'h0000498F : data <= 8'b00000000 ;
			15'h00004990 : data <= 8'b00000000 ;
			15'h00004991 : data <= 8'b00000000 ;
			15'h00004992 : data <= 8'b00000000 ;
			15'h00004993 : data <= 8'b00000000 ;
			15'h00004994 : data <= 8'b00000000 ;
			15'h00004995 : data <= 8'b00000000 ;
			15'h00004996 : data <= 8'b00000000 ;
			15'h00004997 : data <= 8'b00000000 ;
			15'h00004998 : data <= 8'b00000000 ;
			15'h00004999 : data <= 8'b00000000 ;
			15'h0000499A : data <= 8'b00000000 ;
			15'h0000499B : data <= 8'b00000000 ;
			15'h0000499C : data <= 8'b00000000 ;
			15'h0000499D : data <= 8'b00000000 ;
			15'h0000499E : data <= 8'b00000000 ;
			15'h0000499F : data <= 8'b00000000 ;
			15'h000049A0 : data <= 8'b00000000 ;
			15'h000049A1 : data <= 8'b00000000 ;
			15'h000049A2 : data <= 8'b00000000 ;
			15'h000049A3 : data <= 8'b00000000 ;
			15'h000049A4 : data <= 8'b00000000 ;
			15'h000049A5 : data <= 8'b00000000 ;
			15'h000049A6 : data <= 8'b00000000 ;
			15'h000049A7 : data <= 8'b00000000 ;
			15'h000049A8 : data <= 8'b00000000 ;
			15'h000049A9 : data <= 8'b00000000 ;
			15'h000049AA : data <= 8'b00000000 ;
			15'h000049AB : data <= 8'b00000000 ;
			15'h000049AC : data <= 8'b00000000 ;
			15'h000049AD : data <= 8'b00000000 ;
			15'h000049AE : data <= 8'b00000000 ;
			15'h000049AF : data <= 8'b00000000 ;
			15'h000049B0 : data <= 8'b00000000 ;
			15'h000049B1 : data <= 8'b00000000 ;
			15'h000049B2 : data <= 8'b00000000 ;
			15'h000049B3 : data <= 8'b00000000 ;
			15'h000049B4 : data <= 8'b00000000 ;
			15'h000049B5 : data <= 8'b00000000 ;
			15'h000049B6 : data <= 8'b00000000 ;
			15'h000049B7 : data <= 8'b00000000 ;
			15'h000049B8 : data <= 8'b00000000 ;
			15'h000049B9 : data <= 8'b00000000 ;
			15'h000049BA : data <= 8'b00000000 ;
			15'h000049BB : data <= 8'b00000000 ;
			15'h000049BC : data <= 8'b00000000 ;
			15'h000049BD : data <= 8'b00000000 ;
			15'h000049BE : data <= 8'b00000000 ;
			15'h000049BF : data <= 8'b00000000 ;
			15'h000049C0 : data <= 8'b00000000 ;
			15'h000049C1 : data <= 8'b00000000 ;
			15'h000049C2 : data <= 8'b00000000 ;
			15'h000049C3 : data <= 8'b00000000 ;
			15'h000049C4 : data <= 8'b00000000 ;
			15'h000049C5 : data <= 8'b00000000 ;
			15'h000049C6 : data <= 8'b00000000 ;
			15'h000049C7 : data <= 8'b00000000 ;
			15'h000049C8 : data <= 8'b00000000 ;
			15'h000049C9 : data <= 8'b00000000 ;
			15'h000049CA : data <= 8'b00000000 ;
			15'h000049CB : data <= 8'b00000000 ;
			15'h000049CC : data <= 8'b00000000 ;
			15'h000049CD : data <= 8'b00000000 ;
			15'h000049CE : data <= 8'b00000000 ;
			15'h000049CF : data <= 8'b00000000 ;
			15'h000049D0 : data <= 8'b00000000 ;
			15'h000049D1 : data <= 8'b00000000 ;
			15'h000049D2 : data <= 8'b00000000 ;
			15'h000049D3 : data <= 8'b00000000 ;
			15'h000049D4 : data <= 8'b00000000 ;
			15'h000049D5 : data <= 8'b00000000 ;
			15'h000049D6 : data <= 8'b00000000 ;
			15'h000049D7 : data <= 8'b00000000 ;
			15'h000049D8 : data <= 8'b00000000 ;
			15'h000049D9 : data <= 8'b00000000 ;
			15'h000049DA : data <= 8'b00000000 ;
			15'h000049DB : data <= 8'b00000000 ;
			15'h000049DC : data <= 8'b00000000 ;
			15'h000049DD : data <= 8'b00000000 ;
			15'h000049DE : data <= 8'b00000000 ;
			15'h000049DF : data <= 8'b00000000 ;
			15'h000049E0 : data <= 8'b00000000 ;
			15'h000049E1 : data <= 8'b00000000 ;
			15'h000049E2 : data <= 8'b00000000 ;
			15'h000049E3 : data <= 8'b00000000 ;
			15'h000049E4 : data <= 8'b00000000 ;
			15'h000049E5 : data <= 8'b00000000 ;
			15'h000049E6 : data <= 8'b00000000 ;
			15'h000049E7 : data <= 8'b00000000 ;
			15'h000049E8 : data <= 8'b00000000 ;
			15'h000049E9 : data <= 8'b00000000 ;
			15'h000049EA : data <= 8'b00000000 ;
			15'h000049EB : data <= 8'b00000000 ;
			15'h000049EC : data <= 8'b00000000 ;
			15'h000049ED : data <= 8'b00000000 ;
			15'h000049EE : data <= 8'b00000000 ;
			15'h000049EF : data <= 8'b00000000 ;
			15'h000049F0 : data <= 8'b00000000 ;
			15'h000049F1 : data <= 8'b00000000 ;
			15'h000049F2 : data <= 8'b00000000 ;
			15'h000049F3 : data <= 8'b00000000 ;
			15'h000049F4 : data <= 8'b00000000 ;
			15'h000049F5 : data <= 8'b00000000 ;
			15'h000049F6 : data <= 8'b00000000 ;
			15'h000049F7 : data <= 8'b00000000 ;
			15'h000049F8 : data <= 8'b00000000 ;
			15'h000049F9 : data <= 8'b00000000 ;
			15'h000049FA : data <= 8'b00000000 ;
			15'h000049FB : data <= 8'b00000000 ;
			15'h000049FC : data <= 8'b00000000 ;
			15'h000049FD : data <= 8'b00000000 ;
			15'h000049FE : data <= 8'b00000000 ;
			15'h000049FF : data <= 8'b00000000 ;
			15'h00004A00 : data <= 8'b00000000 ;
			15'h00004A01 : data <= 8'b00000000 ;
			15'h00004A02 : data <= 8'b00000000 ;
			15'h00004A03 : data <= 8'b00000000 ;
			15'h00004A04 : data <= 8'b00000000 ;
			15'h00004A05 : data <= 8'b00000000 ;
			15'h00004A06 : data <= 8'b00000000 ;
			15'h00004A07 : data <= 8'b00000000 ;
			15'h00004A08 : data <= 8'b00000000 ;
			15'h00004A09 : data <= 8'b00000000 ;
			15'h00004A0A : data <= 8'b00000000 ;
			15'h00004A0B : data <= 8'b00000000 ;
			15'h00004A0C : data <= 8'b00000000 ;
			15'h00004A0D : data <= 8'b00000000 ;
			15'h00004A0E : data <= 8'b00000000 ;
			15'h00004A0F : data <= 8'b00000000 ;
			15'h00004A10 : data <= 8'b00000000 ;
			15'h00004A11 : data <= 8'b00000000 ;
			15'h00004A12 : data <= 8'b00000000 ;
			15'h00004A13 : data <= 8'b00000000 ;
			15'h00004A14 : data <= 8'b00000000 ;
			15'h00004A15 : data <= 8'b00000000 ;
			15'h00004A16 : data <= 8'b00000000 ;
			15'h00004A17 : data <= 8'b00000000 ;
			15'h00004A18 : data <= 8'b00000000 ;
			15'h00004A19 : data <= 8'b00000000 ;
			15'h00004A1A : data <= 8'b00000000 ;
			15'h00004A1B : data <= 8'b00000000 ;
			15'h00004A1C : data <= 8'b00000000 ;
			15'h00004A1D : data <= 8'b00000000 ;
			15'h00004A1E : data <= 8'b00000000 ;
			15'h00004A1F : data <= 8'b00000000 ;
			15'h00004A20 : data <= 8'b00000000 ;
			15'h00004A21 : data <= 8'b00000000 ;
			15'h00004A22 : data <= 8'b00000000 ;
			15'h00004A23 : data <= 8'b00000000 ;
			15'h00004A24 : data <= 8'b00000000 ;
			15'h00004A25 : data <= 8'b00000000 ;
			15'h00004A26 : data <= 8'b00000000 ;
			15'h00004A27 : data <= 8'b00000000 ;
			15'h00004A28 : data <= 8'b00000000 ;
			15'h00004A29 : data <= 8'b00000000 ;
			15'h00004A2A : data <= 8'b00000000 ;
			15'h00004A2B : data <= 8'b00000000 ;
			15'h00004A2C : data <= 8'b00000000 ;
			15'h00004A2D : data <= 8'b00000000 ;
			15'h00004A2E : data <= 8'b00000000 ;
			15'h00004A2F : data <= 8'b00000000 ;
			15'h00004A30 : data <= 8'b00000000 ;
			15'h00004A31 : data <= 8'b00000000 ;
			15'h00004A32 : data <= 8'b00000000 ;
			15'h00004A33 : data <= 8'b00000000 ;
			15'h00004A34 : data <= 8'b00000000 ;
			15'h00004A35 : data <= 8'b00000000 ;
			15'h00004A36 : data <= 8'b00000000 ;
			15'h00004A37 : data <= 8'b00000000 ;
			15'h00004A38 : data <= 8'b00000000 ;
			15'h00004A39 : data <= 8'b00000000 ;
			15'h00004A3A : data <= 8'b00000000 ;
			15'h00004A3B : data <= 8'b00000000 ;
			15'h00004A3C : data <= 8'b00000000 ;
			15'h00004A3D : data <= 8'b00000000 ;
			15'h00004A3E : data <= 8'b00000000 ;
			15'h00004A3F : data <= 8'b00000000 ;
			15'h00004A40 : data <= 8'b00000000 ;
			15'h00004A41 : data <= 8'b00000000 ;
			15'h00004A42 : data <= 8'b00000000 ;
			15'h00004A43 : data <= 8'b00000000 ;
			15'h00004A44 : data <= 8'b00000000 ;
			15'h00004A45 : data <= 8'b00000000 ;
			15'h00004A46 : data <= 8'b00000000 ;
			15'h00004A47 : data <= 8'b00000000 ;
			15'h00004A48 : data <= 8'b00000000 ;
			15'h00004A49 : data <= 8'b00000000 ;
			15'h00004A4A : data <= 8'b00000000 ;
			15'h00004A4B : data <= 8'b00000000 ;
			15'h00004A4C : data <= 8'b00000000 ;
			15'h00004A4D : data <= 8'b00000000 ;
			15'h00004A4E : data <= 8'b00000000 ;
			15'h00004A4F : data <= 8'b00000000 ;
			15'h00004A50 : data <= 8'b00000000 ;
			15'h00004A51 : data <= 8'b00000000 ;
			15'h00004A52 : data <= 8'b00000000 ;
			15'h00004A53 : data <= 8'b00000000 ;
			15'h00004A54 : data <= 8'b00000000 ;
			15'h00004A55 : data <= 8'b00000000 ;
			15'h00004A56 : data <= 8'b00000000 ;
			15'h00004A57 : data <= 8'b00000000 ;
			15'h00004A58 : data <= 8'b00000000 ;
			15'h00004A59 : data <= 8'b00000000 ;
			15'h00004A5A : data <= 8'b00000000 ;
			15'h00004A5B : data <= 8'b00000000 ;
			15'h00004A5C : data <= 8'b00000000 ;
			15'h00004A5D : data <= 8'b00000000 ;
			15'h00004A5E : data <= 8'b00000000 ;
			15'h00004A5F : data <= 8'b00000000 ;
			15'h00004A60 : data <= 8'b00000000 ;
			15'h00004A61 : data <= 8'b00000000 ;
			15'h00004A62 : data <= 8'b00000000 ;
			15'h00004A63 : data <= 8'b00000000 ;
			15'h00004A64 : data <= 8'b00000000 ;
			15'h00004A65 : data <= 8'b00000000 ;
			15'h00004A66 : data <= 8'b00000000 ;
			15'h00004A67 : data <= 8'b00000000 ;
			15'h00004A68 : data <= 8'b00000000 ;
			15'h00004A69 : data <= 8'b00000000 ;
			15'h00004A6A : data <= 8'b00000000 ;
			15'h00004A6B : data <= 8'b00000000 ;
			15'h00004A6C : data <= 8'b00000000 ;
			15'h00004A6D : data <= 8'b00000000 ;
			15'h00004A6E : data <= 8'b00000000 ;
			15'h00004A6F : data <= 8'b00000000 ;
			15'h00004A70 : data <= 8'b00000000 ;
			15'h00004A71 : data <= 8'b00000000 ;
			15'h00004A72 : data <= 8'b00000000 ;
			15'h00004A73 : data <= 8'b00000000 ;
			15'h00004A74 : data <= 8'b00000000 ;
			15'h00004A75 : data <= 8'b00000000 ;
			15'h00004A76 : data <= 8'b00000000 ;
			15'h00004A77 : data <= 8'b00000000 ;
			15'h00004A78 : data <= 8'b00000000 ;
			15'h00004A79 : data <= 8'b00000000 ;
			15'h00004A7A : data <= 8'b00000000 ;
			15'h00004A7B : data <= 8'b00000000 ;
			15'h00004A7C : data <= 8'b00000000 ;
			15'h00004A7D : data <= 8'b00000000 ;
			15'h00004A7E : data <= 8'b00000000 ;
			15'h00004A7F : data <= 8'b00000000 ;
			15'h00004A80 : data <= 8'b00000000 ;
			15'h00004A81 : data <= 8'b00000000 ;
			15'h00004A82 : data <= 8'b00000000 ;
			15'h00004A83 : data <= 8'b00000000 ;
			15'h00004A84 : data <= 8'b00000000 ;
			15'h00004A85 : data <= 8'b00000000 ;
			15'h00004A86 : data <= 8'b00000000 ;
			15'h00004A87 : data <= 8'b00000000 ;
			15'h00004A88 : data <= 8'b00000000 ;
			15'h00004A89 : data <= 8'b00000000 ;
			15'h00004A8A : data <= 8'b00000000 ;
			15'h00004A8B : data <= 8'b00000000 ;
			15'h00004A8C : data <= 8'b00000000 ;
			15'h00004A8D : data <= 8'b00000000 ;
			15'h00004A8E : data <= 8'b00000000 ;
			15'h00004A8F : data <= 8'b00000000 ;
			15'h00004A90 : data <= 8'b00000000 ;
			15'h00004A91 : data <= 8'b00000000 ;
			15'h00004A92 : data <= 8'b00000000 ;
			15'h00004A93 : data <= 8'b00000000 ;
			15'h00004A94 : data <= 8'b00000000 ;
			15'h00004A95 : data <= 8'b00000000 ;
			15'h00004A96 : data <= 8'b00000000 ;
			15'h00004A97 : data <= 8'b00000000 ;
			15'h00004A98 : data <= 8'b00000000 ;
			15'h00004A99 : data <= 8'b00000000 ;
			15'h00004A9A : data <= 8'b00000000 ;
			15'h00004A9B : data <= 8'b00000000 ;
			15'h00004A9C : data <= 8'b00000000 ;
			15'h00004A9D : data <= 8'b00000000 ;
			15'h00004A9E : data <= 8'b00000000 ;
			15'h00004A9F : data <= 8'b00000000 ;
			15'h00004AA0 : data <= 8'b00000000 ;
			15'h00004AA1 : data <= 8'b00000000 ;
			15'h00004AA2 : data <= 8'b00000000 ;
			15'h00004AA3 : data <= 8'b00000000 ;
			15'h00004AA4 : data <= 8'b00000000 ;
			15'h00004AA5 : data <= 8'b00000000 ;
			15'h00004AA6 : data <= 8'b00000000 ;
			15'h00004AA7 : data <= 8'b00000000 ;
			15'h00004AA8 : data <= 8'b00000000 ;
			15'h00004AA9 : data <= 8'b00000000 ;
			15'h00004AAA : data <= 8'b00000000 ;
			15'h00004AAB : data <= 8'b00000000 ;
			15'h00004AAC : data <= 8'b00000000 ;
			15'h00004AAD : data <= 8'b00000000 ;
			15'h00004AAE : data <= 8'b00000000 ;
			15'h00004AAF : data <= 8'b00000000 ;
			15'h00004AB0 : data <= 8'b00000000 ;
			15'h00004AB1 : data <= 8'b00000000 ;
			15'h00004AB2 : data <= 8'b00000000 ;
			15'h00004AB3 : data <= 8'b00000000 ;
			15'h00004AB4 : data <= 8'b00000000 ;
			15'h00004AB5 : data <= 8'b00000000 ;
			15'h00004AB6 : data <= 8'b00000000 ;
			15'h00004AB7 : data <= 8'b00000000 ;
			15'h00004AB8 : data <= 8'b00000000 ;
			15'h00004AB9 : data <= 8'b00000000 ;
			15'h00004ABA : data <= 8'b00000000 ;
			15'h00004ABB : data <= 8'b00000000 ;
			15'h00004ABC : data <= 8'b00000000 ;
			15'h00004ABD : data <= 8'b00000000 ;
			15'h00004ABE : data <= 8'b00000000 ;
			15'h00004ABF : data <= 8'b00000000 ;
			15'h00004AC0 : data <= 8'b00000000 ;
			15'h00004AC1 : data <= 8'b00000000 ;
			15'h00004AC2 : data <= 8'b00000000 ;
			15'h00004AC3 : data <= 8'b00000000 ;
			15'h00004AC4 : data <= 8'b00000000 ;
			15'h00004AC5 : data <= 8'b00000000 ;
			15'h00004AC6 : data <= 8'b00000000 ;
			15'h00004AC7 : data <= 8'b00000000 ;
			15'h00004AC8 : data <= 8'b00000000 ;
			15'h00004AC9 : data <= 8'b00000000 ;
			15'h00004ACA : data <= 8'b00000000 ;
			15'h00004ACB : data <= 8'b00000000 ;
			15'h00004ACC : data <= 8'b00000000 ;
			15'h00004ACD : data <= 8'b00000000 ;
			15'h00004ACE : data <= 8'b00000000 ;
			15'h00004ACF : data <= 8'b00000000 ;
			15'h00004AD0 : data <= 8'b00000000 ;
			15'h00004AD1 : data <= 8'b00000000 ;
			15'h00004AD2 : data <= 8'b00000000 ;
			15'h00004AD3 : data <= 8'b00000000 ;
			15'h00004AD4 : data <= 8'b00000000 ;
			15'h00004AD5 : data <= 8'b00000000 ;
			15'h00004AD6 : data <= 8'b00000000 ;
			15'h00004AD7 : data <= 8'b00000000 ;
			15'h00004AD8 : data <= 8'b00000000 ;
			15'h00004AD9 : data <= 8'b00000000 ;
			15'h00004ADA : data <= 8'b00000000 ;
			15'h00004ADB : data <= 8'b00000000 ;
			15'h00004ADC : data <= 8'b00000000 ;
			15'h00004ADD : data <= 8'b00000000 ;
			15'h00004ADE : data <= 8'b00000000 ;
			15'h00004ADF : data <= 8'b00000000 ;
			15'h00004AE0 : data <= 8'b00000000 ;
			15'h00004AE1 : data <= 8'b00000000 ;
			15'h00004AE2 : data <= 8'b00000000 ;
			15'h00004AE3 : data <= 8'b00000000 ;
			15'h00004AE4 : data <= 8'b00000000 ;
			15'h00004AE5 : data <= 8'b00000000 ;
			15'h00004AE6 : data <= 8'b00000000 ;
			15'h00004AE7 : data <= 8'b00000000 ;
			15'h00004AE8 : data <= 8'b00000000 ;
			15'h00004AE9 : data <= 8'b00000000 ;
			15'h00004AEA : data <= 8'b00000000 ;
			15'h00004AEB : data <= 8'b00000000 ;
			15'h00004AEC : data <= 8'b00000000 ;
			15'h00004AED : data <= 8'b00000000 ;
			15'h00004AEE : data <= 8'b00000000 ;
			15'h00004AEF : data <= 8'b00000000 ;
			15'h00004AF0 : data <= 8'b00000000 ;
			15'h00004AF1 : data <= 8'b00000000 ;
			15'h00004AF2 : data <= 8'b00000000 ;
			15'h00004AF3 : data <= 8'b00000000 ;
			15'h00004AF4 : data <= 8'b00000000 ;
			15'h00004AF5 : data <= 8'b00000000 ;
			15'h00004AF6 : data <= 8'b00000000 ;
			15'h00004AF7 : data <= 8'b00000000 ;
			15'h00004AF8 : data <= 8'b00000000 ;
			15'h00004AF9 : data <= 8'b00000000 ;
			15'h00004AFA : data <= 8'b00000000 ;
			15'h00004AFB : data <= 8'b00000000 ;
			15'h00004AFC : data <= 8'b00000000 ;
			15'h00004AFD : data <= 8'b00000000 ;
			15'h00004AFE : data <= 8'b00000000 ;
			15'h00004AFF : data <= 8'b00000000 ;
			15'h00004B00 : data <= 8'b00000000 ;
			15'h00004B01 : data <= 8'b00000000 ;
			15'h00004B02 : data <= 8'b00000000 ;
			15'h00004B03 : data <= 8'b00000000 ;
			15'h00004B04 : data <= 8'b00000000 ;
			15'h00004B05 : data <= 8'b00000000 ;
			15'h00004B06 : data <= 8'b00000000 ;
			15'h00004B07 : data <= 8'b00000000 ;
			15'h00004B08 : data <= 8'b00000000 ;
			15'h00004B09 : data <= 8'b00000000 ;
			15'h00004B0A : data <= 8'b00000000 ;
			15'h00004B0B : data <= 8'b00000000 ;
			15'h00004B0C : data <= 8'b00000000 ;
			15'h00004B0D : data <= 8'b00000000 ;
			15'h00004B0E : data <= 8'b00000000 ;
			15'h00004B0F : data <= 8'b00000000 ;
			15'h00004B10 : data <= 8'b00000000 ;
			15'h00004B11 : data <= 8'b00000000 ;
			15'h00004B12 : data <= 8'b00000000 ;
			15'h00004B13 : data <= 8'b00000000 ;
			15'h00004B14 : data <= 8'b00000000 ;
			15'h00004B15 : data <= 8'b00000000 ;
			15'h00004B16 : data <= 8'b00000000 ;
			15'h00004B17 : data <= 8'b00000000 ;
			15'h00004B18 : data <= 8'b00000000 ;
			15'h00004B19 : data <= 8'b00000000 ;
			15'h00004B1A : data <= 8'b00000000 ;
			15'h00004B1B : data <= 8'b00000000 ;
			15'h00004B1C : data <= 8'b00000000 ;
			15'h00004B1D : data <= 8'b00000000 ;
			15'h00004B1E : data <= 8'b00000000 ;
			15'h00004B1F : data <= 8'b00000000 ;
			15'h00004B20 : data <= 8'b00000000 ;
			15'h00004B21 : data <= 8'b00000000 ;
			15'h00004B22 : data <= 8'b00000000 ;
			15'h00004B23 : data <= 8'b00000000 ;
			15'h00004B24 : data <= 8'b00000000 ;
			15'h00004B25 : data <= 8'b00000000 ;
			15'h00004B26 : data <= 8'b00000000 ;
			15'h00004B27 : data <= 8'b00000000 ;
			15'h00004B28 : data <= 8'b00000000 ;
			15'h00004B29 : data <= 8'b00000000 ;
			15'h00004B2A : data <= 8'b00000000 ;
			15'h00004B2B : data <= 8'b00000000 ;
			15'h00004B2C : data <= 8'b00000000 ;
			15'h00004B2D : data <= 8'b00000000 ;
			15'h00004B2E : data <= 8'b00000000 ;
			15'h00004B2F : data <= 8'b00000000 ;
			15'h00004B30 : data <= 8'b00000000 ;
			15'h00004B31 : data <= 8'b00000000 ;
			15'h00004B32 : data <= 8'b00000000 ;
			15'h00004B33 : data <= 8'b00000000 ;
			15'h00004B34 : data <= 8'b00000000 ;
			15'h00004B35 : data <= 8'b00000000 ;
			15'h00004B36 : data <= 8'b00000000 ;
			15'h00004B37 : data <= 8'b00000000 ;
			15'h00004B38 : data <= 8'b00000000 ;
			15'h00004B39 : data <= 8'b00000000 ;
			15'h00004B3A : data <= 8'b00000000 ;
			15'h00004B3B : data <= 8'b00000000 ;
			15'h00004B3C : data <= 8'b00000000 ;
			15'h00004B3D : data <= 8'b00000000 ;
			15'h00004B3E : data <= 8'b00000000 ;
			15'h00004B3F : data <= 8'b00000000 ;
			15'h00004B40 : data <= 8'b00000000 ;
			15'h00004B41 : data <= 8'b00000000 ;
			15'h00004B42 : data <= 8'b00000000 ;
			15'h00004B43 : data <= 8'b00000000 ;
			15'h00004B44 : data <= 8'b00000000 ;
			15'h00004B45 : data <= 8'b00000000 ;
			15'h00004B46 : data <= 8'b00000000 ;
			15'h00004B47 : data <= 8'b00000000 ;
			15'h00004B48 : data <= 8'b00000000 ;
			15'h00004B49 : data <= 8'b00000000 ;
			15'h00004B4A : data <= 8'b00000000 ;
			15'h00004B4B : data <= 8'b00000000 ;
			15'h00004B4C : data <= 8'b00000000 ;
			15'h00004B4D : data <= 8'b00000000 ;
			15'h00004B4E : data <= 8'b00000000 ;
			15'h00004B4F : data <= 8'b00000000 ;
			15'h00004B50 : data <= 8'b00000000 ;
			15'h00004B51 : data <= 8'b00000000 ;
			15'h00004B52 : data <= 8'b00000000 ;
			15'h00004B53 : data <= 8'b00000000 ;
			15'h00004B54 : data <= 8'b00000000 ;
			15'h00004B55 : data <= 8'b00000000 ;
			15'h00004B56 : data <= 8'b00000000 ;
			15'h00004B57 : data <= 8'b00000000 ;
			15'h00004B58 : data <= 8'b00000000 ;
			15'h00004B59 : data <= 8'b00000000 ;
			15'h00004B5A : data <= 8'b00000000 ;
			15'h00004B5B : data <= 8'b00000000 ;
			15'h00004B5C : data <= 8'b00000000 ;
			15'h00004B5D : data <= 8'b00000000 ;
			15'h00004B5E : data <= 8'b00000000 ;
			15'h00004B5F : data <= 8'b00000000 ;
			15'h00004B60 : data <= 8'b00000000 ;
			15'h00004B61 : data <= 8'b00000000 ;
			15'h00004B62 : data <= 8'b00000000 ;
			15'h00004B63 : data <= 8'b00000000 ;
			15'h00004B64 : data <= 8'b00000000 ;
			15'h00004B65 : data <= 8'b00000000 ;
			15'h00004B66 : data <= 8'b00000000 ;
			15'h00004B67 : data <= 8'b00000000 ;
			15'h00004B68 : data <= 8'b00000000 ;
			15'h00004B69 : data <= 8'b00000000 ;
			15'h00004B6A : data <= 8'b00000000 ;
			15'h00004B6B : data <= 8'b00000000 ;
			15'h00004B6C : data <= 8'b00000000 ;
			15'h00004B6D : data <= 8'b00000000 ;
			15'h00004B6E : data <= 8'b00000000 ;
			15'h00004B6F : data <= 8'b00000000 ;
			15'h00004B70 : data <= 8'b00000000 ;
			15'h00004B71 : data <= 8'b00000000 ;
			15'h00004B72 : data <= 8'b00000000 ;
			15'h00004B73 : data <= 8'b00000000 ;
			15'h00004B74 : data <= 8'b00000000 ;
			15'h00004B75 : data <= 8'b00000000 ;
			15'h00004B76 : data <= 8'b00000000 ;
			15'h00004B77 : data <= 8'b00000000 ;
			15'h00004B78 : data <= 8'b00000000 ;
			15'h00004B79 : data <= 8'b00000000 ;
			15'h00004B7A : data <= 8'b00000000 ;
			15'h00004B7B : data <= 8'b00000000 ;
			15'h00004B7C : data <= 8'b00000000 ;
			15'h00004B7D : data <= 8'b00000000 ;
			15'h00004B7E : data <= 8'b00000000 ;
			15'h00004B7F : data <= 8'b00000000 ;
			15'h00004B80 : data <= 8'b00000000 ;
			15'h00004B81 : data <= 8'b00000000 ;
			15'h00004B82 : data <= 8'b00000000 ;
			15'h00004B83 : data <= 8'b00000000 ;
			15'h00004B84 : data <= 8'b00000000 ;
			15'h00004B85 : data <= 8'b00000000 ;
			15'h00004B86 : data <= 8'b00000000 ;
			15'h00004B87 : data <= 8'b00000000 ;
			15'h00004B88 : data <= 8'b00000000 ;
			15'h00004B89 : data <= 8'b00000000 ;
			15'h00004B8A : data <= 8'b00000000 ;
			15'h00004B8B : data <= 8'b00000000 ;
			15'h00004B8C : data <= 8'b00000000 ;
			15'h00004B8D : data <= 8'b00000000 ;
			15'h00004B8E : data <= 8'b00000000 ;
			15'h00004B8F : data <= 8'b00000000 ;
			15'h00004B90 : data <= 8'b00000000 ;
			15'h00004B91 : data <= 8'b00000000 ;
			15'h00004B92 : data <= 8'b00000000 ;
			15'h00004B93 : data <= 8'b00000000 ;
			15'h00004B94 : data <= 8'b00000000 ;
			15'h00004B95 : data <= 8'b00000000 ;
			15'h00004B96 : data <= 8'b00000000 ;
			15'h00004B97 : data <= 8'b00000000 ;
			15'h00004B98 : data <= 8'b00000000 ;
			15'h00004B99 : data <= 8'b00000000 ;
			15'h00004B9A : data <= 8'b00000000 ;
			15'h00004B9B : data <= 8'b00000000 ;
			15'h00004B9C : data <= 8'b00000000 ;
			15'h00004B9D : data <= 8'b00000000 ;
			15'h00004B9E : data <= 8'b00000000 ;
			15'h00004B9F : data <= 8'b00000000 ;
			15'h00004BA0 : data <= 8'b00000000 ;
			15'h00004BA1 : data <= 8'b00000000 ;
			15'h00004BA2 : data <= 8'b00000000 ;
			15'h00004BA3 : data <= 8'b00000000 ;
			15'h00004BA4 : data <= 8'b00000000 ;
			15'h00004BA5 : data <= 8'b00000000 ;
			15'h00004BA6 : data <= 8'b00000000 ;
			15'h00004BA7 : data <= 8'b00000000 ;
			15'h00004BA8 : data <= 8'b00000000 ;
			15'h00004BA9 : data <= 8'b00000000 ;
			15'h00004BAA : data <= 8'b00000000 ;
			15'h00004BAB : data <= 8'b00000000 ;
			15'h00004BAC : data <= 8'b00000000 ;
			15'h00004BAD : data <= 8'b00000000 ;
			15'h00004BAE : data <= 8'b00000000 ;
			15'h00004BAF : data <= 8'b00000000 ;
			15'h00004BB0 : data <= 8'b00000000 ;
			15'h00004BB1 : data <= 8'b00000000 ;
			15'h00004BB2 : data <= 8'b00000000 ;
			15'h00004BB3 : data <= 8'b00000000 ;
			15'h00004BB4 : data <= 8'b00000000 ;
			15'h00004BB5 : data <= 8'b00000000 ;
			15'h00004BB6 : data <= 8'b00000000 ;
			15'h00004BB7 : data <= 8'b00000000 ;
			15'h00004BB8 : data <= 8'b00000000 ;
			15'h00004BB9 : data <= 8'b00000000 ;
			15'h00004BBA : data <= 8'b00000000 ;
			15'h00004BBB : data <= 8'b00000000 ;
			15'h00004BBC : data <= 8'b00000000 ;
			15'h00004BBD : data <= 8'b00000000 ;
			15'h00004BBE : data <= 8'b00000000 ;
			15'h00004BBF : data <= 8'b00000000 ;
			15'h00004BC0 : data <= 8'b00000000 ;
			15'h00004BC1 : data <= 8'b00000000 ;
			15'h00004BC2 : data <= 8'b00000000 ;
			15'h00004BC3 : data <= 8'b00000000 ;
			15'h00004BC4 : data <= 8'b00000000 ;
			15'h00004BC5 : data <= 8'b00000000 ;
			15'h00004BC6 : data <= 8'b00000000 ;
			15'h00004BC7 : data <= 8'b00000000 ;
			15'h00004BC8 : data <= 8'b00000000 ;
			15'h00004BC9 : data <= 8'b00000000 ;
			15'h00004BCA : data <= 8'b00000000 ;
			15'h00004BCB : data <= 8'b00000000 ;
			15'h00004BCC : data <= 8'b00000000 ;
			15'h00004BCD : data <= 8'b00000000 ;
			15'h00004BCE : data <= 8'b00000000 ;
			15'h00004BCF : data <= 8'b00000000 ;
			15'h00004BD0 : data <= 8'b00000000 ;
			15'h00004BD1 : data <= 8'b00000000 ;
			15'h00004BD2 : data <= 8'b00000000 ;
			15'h00004BD3 : data <= 8'b00000000 ;
			15'h00004BD4 : data <= 8'b00000000 ;
			15'h00004BD5 : data <= 8'b00000000 ;
			15'h00004BD6 : data <= 8'b00000000 ;
			15'h00004BD7 : data <= 8'b00000000 ;
			15'h00004BD8 : data <= 8'b00000000 ;
			15'h00004BD9 : data <= 8'b00000000 ;
			15'h00004BDA : data <= 8'b00000000 ;
			15'h00004BDB : data <= 8'b00000000 ;
			15'h00004BDC : data <= 8'b00000000 ;
			15'h00004BDD : data <= 8'b00000000 ;
			15'h00004BDE : data <= 8'b00000000 ;
			15'h00004BDF : data <= 8'b00000000 ;
			15'h00004BE0 : data <= 8'b00000000 ;
			15'h00004BE1 : data <= 8'b00000000 ;
			15'h00004BE2 : data <= 8'b00000000 ;
			15'h00004BE3 : data <= 8'b00000000 ;
			15'h00004BE4 : data <= 8'b00000000 ;
			15'h00004BE5 : data <= 8'b00000000 ;
			15'h00004BE6 : data <= 8'b00000000 ;
			15'h00004BE7 : data <= 8'b00000000 ;
			15'h00004BE8 : data <= 8'b00000000 ;
			15'h00004BE9 : data <= 8'b00000000 ;
			15'h00004BEA : data <= 8'b00000000 ;
			15'h00004BEB : data <= 8'b00000000 ;
			15'h00004BEC : data <= 8'b00000000 ;
			15'h00004BED : data <= 8'b00000000 ;
			15'h00004BEE : data <= 8'b00000000 ;
			15'h00004BEF : data <= 8'b00000000 ;
			15'h00004BF0 : data <= 8'b00000000 ;
			15'h00004BF1 : data <= 8'b00000000 ;
			15'h00004BF2 : data <= 8'b00000000 ;
			15'h00004BF3 : data <= 8'b00000000 ;
			15'h00004BF4 : data <= 8'b00000000 ;
			15'h00004BF5 : data <= 8'b00000000 ;
			15'h00004BF6 : data <= 8'b00000000 ;
			15'h00004BF7 : data <= 8'b00000000 ;
			15'h00004BF8 : data <= 8'b00000000 ;
			15'h00004BF9 : data <= 8'b00000000 ;
			15'h00004BFA : data <= 8'b00000000 ;
			15'h00004BFB : data <= 8'b00000000 ;
			15'h00004BFC : data <= 8'b00000000 ;
			15'h00004BFD : data <= 8'b00000000 ;
			15'h00004BFE : data <= 8'b00000000 ;
			15'h00004BFF : data <= 8'b00000000 ;
			15'h00004C00 : data <= 8'b00000000 ;
			15'h00004C01 : data <= 8'b00000000 ;
			15'h00004C02 : data <= 8'b00000000 ;
			15'h00004C03 : data <= 8'b00000000 ;
			15'h00004C04 : data <= 8'b00000000 ;
			15'h00004C05 : data <= 8'b00000000 ;
			15'h00004C06 : data <= 8'b00000000 ;
			15'h00004C07 : data <= 8'b00000000 ;
			15'h00004C08 : data <= 8'b00000000 ;
			15'h00004C09 : data <= 8'b00000000 ;
			15'h00004C0A : data <= 8'b00000000 ;
			15'h00004C0B : data <= 8'b00000000 ;
			15'h00004C0C : data <= 8'b00000000 ;
			15'h00004C0D : data <= 8'b00000000 ;
			15'h00004C0E : data <= 8'b00000000 ;
			15'h00004C0F : data <= 8'b00000000 ;
			15'h00004C10 : data <= 8'b00000000 ;
			15'h00004C11 : data <= 8'b00000000 ;
			15'h00004C12 : data <= 8'b00000000 ;
			15'h00004C13 : data <= 8'b00000000 ;
			15'h00004C14 : data <= 8'b00000000 ;
			15'h00004C15 : data <= 8'b00000000 ;
			15'h00004C16 : data <= 8'b00000000 ;
			15'h00004C17 : data <= 8'b00000000 ;
			15'h00004C18 : data <= 8'b00000000 ;
			15'h00004C19 : data <= 8'b00000000 ;
			15'h00004C1A : data <= 8'b00000000 ;
			15'h00004C1B : data <= 8'b00000000 ;
			15'h00004C1C : data <= 8'b00000000 ;
			15'h00004C1D : data <= 8'b00000000 ;
			15'h00004C1E : data <= 8'b00000000 ;
			15'h00004C1F : data <= 8'b00000000 ;
			15'h00004C20 : data <= 8'b00000000 ;
			15'h00004C21 : data <= 8'b00000000 ;
			15'h00004C22 : data <= 8'b00000000 ;
			15'h00004C23 : data <= 8'b00000000 ;
			15'h00004C24 : data <= 8'b00000000 ;
			15'h00004C25 : data <= 8'b00000000 ;
			15'h00004C26 : data <= 8'b00000000 ;
			15'h00004C27 : data <= 8'b00000000 ;
			15'h00004C28 : data <= 8'b00000000 ;
			15'h00004C29 : data <= 8'b00000000 ;
			15'h00004C2A : data <= 8'b00000000 ;
			15'h00004C2B : data <= 8'b00000000 ;
			15'h00004C2C : data <= 8'b00000000 ;
			15'h00004C2D : data <= 8'b00000000 ;
			15'h00004C2E : data <= 8'b00000000 ;
			15'h00004C2F : data <= 8'b00000000 ;
			15'h00004C30 : data <= 8'b00000000 ;
			15'h00004C31 : data <= 8'b00000000 ;
			15'h00004C32 : data <= 8'b00000000 ;
			15'h00004C33 : data <= 8'b00000000 ;
			15'h00004C34 : data <= 8'b00000000 ;
			15'h00004C35 : data <= 8'b00000000 ;
			15'h00004C36 : data <= 8'b00000000 ;
			15'h00004C37 : data <= 8'b00000000 ;
			15'h00004C38 : data <= 8'b00000000 ;
			15'h00004C39 : data <= 8'b00000000 ;
			15'h00004C3A : data <= 8'b00000000 ;
			15'h00004C3B : data <= 8'b00000000 ;
			15'h00004C3C : data <= 8'b00000000 ;
			15'h00004C3D : data <= 8'b00000000 ;
			15'h00004C3E : data <= 8'b00000000 ;
			15'h00004C3F : data <= 8'b00000000 ;
			15'h00004C40 : data <= 8'b00000000 ;
			15'h00004C41 : data <= 8'b00000000 ;
			15'h00004C42 : data <= 8'b00000000 ;
			15'h00004C43 : data <= 8'b00000000 ;
			15'h00004C44 : data <= 8'b00000000 ;
			15'h00004C45 : data <= 8'b00000000 ;
			15'h00004C46 : data <= 8'b00000000 ;
			15'h00004C47 : data <= 8'b00000000 ;
			15'h00004C48 : data <= 8'b00000000 ;
			15'h00004C49 : data <= 8'b00000000 ;
			15'h00004C4A : data <= 8'b00000000 ;
			15'h00004C4B : data <= 8'b00000000 ;
			15'h00004C4C : data <= 8'b00000000 ;
			15'h00004C4D : data <= 8'b00000000 ;
			15'h00004C4E : data <= 8'b00000000 ;
			15'h00004C4F : data <= 8'b00000000 ;
			15'h00004C50 : data <= 8'b00000000 ;
			15'h00004C51 : data <= 8'b00000000 ;
			15'h00004C52 : data <= 8'b00000000 ;
			15'h00004C53 : data <= 8'b00000000 ;
			15'h00004C54 : data <= 8'b00000000 ;
			15'h00004C55 : data <= 8'b00000000 ;
			15'h00004C56 : data <= 8'b00000000 ;
			15'h00004C57 : data <= 8'b00000000 ;
			15'h00004C58 : data <= 8'b00000000 ;
			15'h00004C59 : data <= 8'b00000000 ;
			15'h00004C5A : data <= 8'b00000000 ;
			15'h00004C5B : data <= 8'b00000000 ;
			15'h00004C5C : data <= 8'b00000000 ;
			15'h00004C5D : data <= 8'b00000000 ;
			15'h00004C5E : data <= 8'b00000000 ;
			15'h00004C5F : data <= 8'b00000000 ;
			15'h00004C60 : data <= 8'b00000000 ;
			15'h00004C61 : data <= 8'b00000000 ;
			15'h00004C62 : data <= 8'b00000000 ;
			15'h00004C63 : data <= 8'b00000000 ;
			15'h00004C64 : data <= 8'b00000000 ;
			15'h00004C65 : data <= 8'b00000000 ;
			15'h00004C66 : data <= 8'b00000000 ;
			15'h00004C67 : data <= 8'b00000000 ;
			15'h00004C68 : data <= 8'b00000000 ;
			15'h00004C69 : data <= 8'b00000000 ;
			15'h00004C6A : data <= 8'b00000000 ;
			15'h00004C6B : data <= 8'b00000000 ;
			15'h00004C6C : data <= 8'b00000000 ;
			15'h00004C6D : data <= 8'b00000000 ;
			15'h00004C6E : data <= 8'b00000000 ;
			15'h00004C6F : data <= 8'b00000000 ;
			15'h00004C70 : data <= 8'b00000000 ;
			15'h00004C71 : data <= 8'b00000000 ;
			15'h00004C72 : data <= 8'b00000000 ;
			15'h00004C73 : data <= 8'b00000000 ;
			15'h00004C74 : data <= 8'b00000000 ;
			15'h00004C75 : data <= 8'b00000000 ;
			15'h00004C76 : data <= 8'b00000000 ;
			15'h00004C77 : data <= 8'b00000000 ;
			15'h00004C78 : data <= 8'b00000000 ;
			15'h00004C79 : data <= 8'b00000000 ;
			15'h00004C7A : data <= 8'b00000000 ;
			15'h00004C7B : data <= 8'b00000000 ;
			15'h00004C7C : data <= 8'b00000000 ;
			15'h00004C7D : data <= 8'b00000000 ;
			15'h00004C7E : data <= 8'b00000000 ;
			15'h00004C7F : data <= 8'b00000000 ;
			15'h00004C80 : data <= 8'b00000000 ;
			15'h00004C81 : data <= 8'b00000000 ;
			15'h00004C82 : data <= 8'b00000000 ;
			15'h00004C83 : data <= 8'b00000000 ;
			15'h00004C84 : data <= 8'b00000000 ;
			15'h00004C85 : data <= 8'b00000000 ;
			15'h00004C86 : data <= 8'b00000000 ;
			15'h00004C87 : data <= 8'b00000000 ;
			15'h00004C88 : data <= 8'b00000000 ;
			15'h00004C89 : data <= 8'b00000000 ;
			15'h00004C8A : data <= 8'b00000000 ;
			15'h00004C8B : data <= 8'b00000000 ;
			15'h00004C8C : data <= 8'b00000000 ;
			15'h00004C8D : data <= 8'b00000000 ;
			15'h00004C8E : data <= 8'b00000000 ;
			15'h00004C8F : data <= 8'b00000000 ;
			15'h00004C90 : data <= 8'b00000000 ;
			15'h00004C91 : data <= 8'b00000000 ;
			15'h00004C92 : data <= 8'b00000000 ;
			15'h00004C93 : data <= 8'b00000000 ;
			15'h00004C94 : data <= 8'b00000000 ;
			15'h00004C95 : data <= 8'b00000000 ;
			15'h00004C96 : data <= 8'b00000000 ;
			15'h00004C97 : data <= 8'b00000000 ;
			15'h00004C98 : data <= 8'b00000000 ;
			15'h00004C99 : data <= 8'b00000000 ;
			15'h00004C9A : data <= 8'b00000000 ;
			15'h00004C9B : data <= 8'b00000000 ;
			15'h00004C9C : data <= 8'b00000000 ;
			15'h00004C9D : data <= 8'b00000000 ;
			15'h00004C9E : data <= 8'b00000000 ;
			15'h00004C9F : data <= 8'b00000000 ;
			15'h00004CA0 : data <= 8'b00000000 ;
			15'h00004CA1 : data <= 8'b00000000 ;
			15'h00004CA2 : data <= 8'b00000000 ;
			15'h00004CA3 : data <= 8'b00000000 ;
			15'h00004CA4 : data <= 8'b00000000 ;
			15'h00004CA5 : data <= 8'b00000000 ;
			15'h00004CA6 : data <= 8'b00000000 ;
			15'h00004CA7 : data <= 8'b00000000 ;
			15'h00004CA8 : data <= 8'b00000000 ;
			15'h00004CA9 : data <= 8'b00000000 ;
			15'h00004CAA : data <= 8'b00000000 ;
			15'h00004CAB : data <= 8'b00000000 ;
			15'h00004CAC : data <= 8'b00000000 ;
			15'h00004CAD : data <= 8'b00000000 ;
			15'h00004CAE : data <= 8'b00000000 ;
			15'h00004CAF : data <= 8'b00000000 ;
			15'h00004CB0 : data <= 8'b00000000 ;
			15'h00004CB1 : data <= 8'b00000000 ;
			15'h00004CB2 : data <= 8'b00000000 ;
			15'h00004CB3 : data <= 8'b00000000 ;
			15'h00004CB4 : data <= 8'b00000000 ;
			15'h00004CB5 : data <= 8'b00000000 ;
			15'h00004CB6 : data <= 8'b00000000 ;
			15'h00004CB7 : data <= 8'b00000000 ;
			15'h00004CB8 : data <= 8'b00000000 ;
			15'h00004CB9 : data <= 8'b00000000 ;
			15'h00004CBA : data <= 8'b00000000 ;
			15'h00004CBB : data <= 8'b00000000 ;
			15'h00004CBC : data <= 8'b00000000 ;
			15'h00004CBD : data <= 8'b00000000 ;
			15'h00004CBE : data <= 8'b00000000 ;
			15'h00004CBF : data <= 8'b00000000 ;
			15'h00004CC0 : data <= 8'b00000000 ;
			15'h00004CC1 : data <= 8'b00000000 ;
			15'h00004CC2 : data <= 8'b00000000 ;
			15'h00004CC3 : data <= 8'b00000000 ;
			15'h00004CC4 : data <= 8'b00000000 ;
			15'h00004CC5 : data <= 8'b00000000 ;
			15'h00004CC6 : data <= 8'b00000000 ;
			15'h00004CC7 : data <= 8'b00000000 ;
			15'h00004CC8 : data <= 8'b00000000 ;
			15'h00004CC9 : data <= 8'b00000000 ;
			15'h00004CCA : data <= 8'b00000000 ;
			15'h00004CCB : data <= 8'b00000000 ;
			15'h00004CCC : data <= 8'b00000000 ;
			15'h00004CCD : data <= 8'b00000000 ;
			15'h00004CCE : data <= 8'b00000000 ;
			15'h00004CCF : data <= 8'b00000000 ;
			15'h00004CD0 : data <= 8'b00000000 ;
			15'h00004CD1 : data <= 8'b00000000 ;
			15'h00004CD2 : data <= 8'b00000000 ;
			15'h00004CD3 : data <= 8'b00000000 ;
			15'h00004CD4 : data <= 8'b00000000 ;
			15'h00004CD5 : data <= 8'b00000000 ;
			15'h00004CD6 : data <= 8'b00000000 ;
			15'h00004CD7 : data <= 8'b00000000 ;
			15'h00004CD8 : data <= 8'b00000000 ;
			15'h00004CD9 : data <= 8'b00000000 ;
			15'h00004CDA : data <= 8'b00000000 ;
			15'h00004CDB : data <= 8'b00000000 ;
			15'h00004CDC : data <= 8'b00000000 ;
			15'h00004CDD : data <= 8'b00000000 ;
			15'h00004CDE : data <= 8'b00000000 ;
			15'h00004CDF : data <= 8'b00000000 ;
			15'h00004CE0 : data <= 8'b00000000 ;
			15'h00004CE1 : data <= 8'b00000000 ;
			15'h00004CE2 : data <= 8'b00000000 ;
			15'h00004CE3 : data <= 8'b00000000 ;
			15'h00004CE4 : data <= 8'b00000000 ;
			15'h00004CE5 : data <= 8'b00000000 ;
			15'h00004CE6 : data <= 8'b00000000 ;
			15'h00004CE7 : data <= 8'b00000000 ;
			15'h00004CE8 : data <= 8'b00000000 ;
			15'h00004CE9 : data <= 8'b00000000 ;
			15'h00004CEA : data <= 8'b00000000 ;
			15'h00004CEB : data <= 8'b00000000 ;
			15'h00004CEC : data <= 8'b00000000 ;
			15'h00004CED : data <= 8'b00000000 ;
			15'h00004CEE : data <= 8'b00000000 ;
			15'h00004CEF : data <= 8'b00000000 ;
			15'h00004CF0 : data <= 8'b00000000 ;
			15'h00004CF1 : data <= 8'b00000000 ;
			15'h00004CF2 : data <= 8'b00000000 ;
			15'h00004CF3 : data <= 8'b00000000 ;
			15'h00004CF4 : data <= 8'b00000000 ;
			15'h00004CF5 : data <= 8'b00000000 ;
			15'h00004CF6 : data <= 8'b00000000 ;
			15'h00004CF7 : data <= 8'b00000000 ;
			15'h00004CF8 : data <= 8'b00000000 ;
			15'h00004CF9 : data <= 8'b00000000 ;
			15'h00004CFA : data <= 8'b00000000 ;
			15'h00004CFB : data <= 8'b00000000 ;
			15'h00004CFC : data <= 8'b00000000 ;
			15'h00004CFD : data <= 8'b00000000 ;
			15'h00004CFE : data <= 8'b00000000 ;
			15'h00004CFF : data <= 8'b00000000 ;
			15'h00004D00 : data <= 8'b00000000 ;
			15'h00004D01 : data <= 8'b00000000 ;
			15'h00004D02 : data <= 8'b00000000 ;
			15'h00004D03 : data <= 8'b00000000 ;
			15'h00004D04 : data <= 8'b00000000 ;
			15'h00004D05 : data <= 8'b00000000 ;
			15'h00004D06 : data <= 8'b00000000 ;
			15'h00004D07 : data <= 8'b00000000 ;
			15'h00004D08 : data <= 8'b00000000 ;
			15'h00004D09 : data <= 8'b00000000 ;
			15'h00004D0A : data <= 8'b00000000 ;
			15'h00004D0B : data <= 8'b00000000 ;
			15'h00004D0C : data <= 8'b00000000 ;
			15'h00004D0D : data <= 8'b00000000 ;
			15'h00004D0E : data <= 8'b00000000 ;
			15'h00004D0F : data <= 8'b00000000 ;
			15'h00004D10 : data <= 8'b00000000 ;
			15'h00004D11 : data <= 8'b00000000 ;
			15'h00004D12 : data <= 8'b00000000 ;
			15'h00004D13 : data <= 8'b00000000 ;
			15'h00004D14 : data <= 8'b00000000 ;
			15'h00004D15 : data <= 8'b00000000 ;
			15'h00004D16 : data <= 8'b00000000 ;
			15'h00004D17 : data <= 8'b00000000 ;
			15'h00004D18 : data <= 8'b00000000 ;
			15'h00004D19 : data <= 8'b00000000 ;
			15'h00004D1A : data <= 8'b00000000 ;
			15'h00004D1B : data <= 8'b00000000 ;
			15'h00004D1C : data <= 8'b00000000 ;
			15'h00004D1D : data <= 8'b00000000 ;
			15'h00004D1E : data <= 8'b00000000 ;
			15'h00004D1F : data <= 8'b00000000 ;
			15'h00004D20 : data <= 8'b00000000 ;
			15'h00004D21 : data <= 8'b00000000 ;
			15'h00004D22 : data <= 8'b00000000 ;
			15'h00004D23 : data <= 8'b00000000 ;
			15'h00004D24 : data <= 8'b00000000 ;
			15'h00004D25 : data <= 8'b00000000 ;
			15'h00004D26 : data <= 8'b00000000 ;
			15'h00004D27 : data <= 8'b00000000 ;
			15'h00004D28 : data <= 8'b00000000 ;
			15'h00004D29 : data <= 8'b00000000 ;
			15'h00004D2A : data <= 8'b00000000 ;
			15'h00004D2B : data <= 8'b00000000 ;
			15'h00004D2C : data <= 8'b00000000 ;
			15'h00004D2D : data <= 8'b00000000 ;
			15'h00004D2E : data <= 8'b00000000 ;
			15'h00004D2F : data <= 8'b00000000 ;
			15'h00004D30 : data <= 8'b00000000 ;
			15'h00004D31 : data <= 8'b00000000 ;
			15'h00004D32 : data <= 8'b00000000 ;
			15'h00004D33 : data <= 8'b00000000 ;
			15'h00004D34 : data <= 8'b00000000 ;
			15'h00004D35 : data <= 8'b00000000 ;
			15'h00004D36 : data <= 8'b00000000 ;
			15'h00004D37 : data <= 8'b00000000 ;
			15'h00004D38 : data <= 8'b00000000 ;
			15'h00004D39 : data <= 8'b00000000 ;
			15'h00004D3A : data <= 8'b00000000 ;
			15'h00004D3B : data <= 8'b00000000 ;
			15'h00004D3C : data <= 8'b00000000 ;
			15'h00004D3D : data <= 8'b00000000 ;
			15'h00004D3E : data <= 8'b00000000 ;
			15'h00004D3F : data <= 8'b00000000 ;
			15'h00004D40 : data <= 8'b00000000 ;
			15'h00004D41 : data <= 8'b00000000 ;
			15'h00004D42 : data <= 8'b00000000 ;
			15'h00004D43 : data <= 8'b00000000 ;
			15'h00004D44 : data <= 8'b00000000 ;
			15'h00004D45 : data <= 8'b00000000 ;
			15'h00004D46 : data <= 8'b00000000 ;
			15'h00004D47 : data <= 8'b00000000 ;
			15'h00004D48 : data <= 8'b00000000 ;
			15'h00004D49 : data <= 8'b00000000 ;
			15'h00004D4A : data <= 8'b00000000 ;
			15'h00004D4B : data <= 8'b00000000 ;
			15'h00004D4C : data <= 8'b00000000 ;
			15'h00004D4D : data <= 8'b00000000 ;
			15'h00004D4E : data <= 8'b00000000 ;
			15'h00004D4F : data <= 8'b00000000 ;
			15'h00004D50 : data <= 8'b00000000 ;
			15'h00004D51 : data <= 8'b00000000 ;
			15'h00004D52 : data <= 8'b00000000 ;
			15'h00004D53 : data <= 8'b00000000 ;
			15'h00004D54 : data <= 8'b00000000 ;
			15'h00004D55 : data <= 8'b00000000 ;
			15'h00004D56 : data <= 8'b00000000 ;
			15'h00004D57 : data <= 8'b00000000 ;
			15'h00004D58 : data <= 8'b00000000 ;
			15'h00004D59 : data <= 8'b00000000 ;
			15'h00004D5A : data <= 8'b00000000 ;
			15'h00004D5B : data <= 8'b00000000 ;
			15'h00004D5C : data <= 8'b00000000 ;
			15'h00004D5D : data <= 8'b00000000 ;
			15'h00004D5E : data <= 8'b00000000 ;
			15'h00004D5F : data <= 8'b00000000 ;
			15'h00004D60 : data <= 8'b00000000 ;
			15'h00004D61 : data <= 8'b00000000 ;
			15'h00004D62 : data <= 8'b00000000 ;
			15'h00004D63 : data <= 8'b00000000 ;
			15'h00004D64 : data <= 8'b00000000 ;
			15'h00004D65 : data <= 8'b00000000 ;
			15'h00004D66 : data <= 8'b00000000 ;
			15'h00004D67 : data <= 8'b00000000 ;
			15'h00004D68 : data <= 8'b00000000 ;
			15'h00004D69 : data <= 8'b00000000 ;
			15'h00004D6A : data <= 8'b00000000 ;
			15'h00004D6B : data <= 8'b00000000 ;
			15'h00004D6C : data <= 8'b00000000 ;
			15'h00004D6D : data <= 8'b00000000 ;
			15'h00004D6E : data <= 8'b00000000 ;
			15'h00004D6F : data <= 8'b00000000 ;
			15'h00004D70 : data <= 8'b00000000 ;
			15'h00004D71 : data <= 8'b00000000 ;
			15'h00004D72 : data <= 8'b00000000 ;
			15'h00004D73 : data <= 8'b00000000 ;
			15'h00004D74 : data <= 8'b00000000 ;
			15'h00004D75 : data <= 8'b00000000 ;
			15'h00004D76 : data <= 8'b00000000 ;
			15'h00004D77 : data <= 8'b00000000 ;
			15'h00004D78 : data <= 8'b00000000 ;
			15'h00004D79 : data <= 8'b00000000 ;
			15'h00004D7A : data <= 8'b00000000 ;
			15'h00004D7B : data <= 8'b00000000 ;
			15'h00004D7C : data <= 8'b00000000 ;
			15'h00004D7D : data <= 8'b00000000 ;
			15'h00004D7E : data <= 8'b00000000 ;
			15'h00004D7F : data <= 8'b00000000 ;
			15'h00004D80 : data <= 8'b00000000 ;
			15'h00004D81 : data <= 8'b00000000 ;
			15'h00004D82 : data <= 8'b00000000 ;
			15'h00004D83 : data <= 8'b00000000 ;
			15'h00004D84 : data <= 8'b00000000 ;
			15'h00004D85 : data <= 8'b00000000 ;
			15'h00004D86 : data <= 8'b00000000 ;
			15'h00004D87 : data <= 8'b00000000 ;
			15'h00004D88 : data <= 8'b00000000 ;
			15'h00004D89 : data <= 8'b00000000 ;
			15'h00004D8A : data <= 8'b00000000 ;
			15'h00004D8B : data <= 8'b00000000 ;
			15'h00004D8C : data <= 8'b00000000 ;
			15'h00004D8D : data <= 8'b00000000 ;
			15'h00004D8E : data <= 8'b00000000 ;
			15'h00004D8F : data <= 8'b00000000 ;
			15'h00004D90 : data <= 8'b00000000 ;
			15'h00004D91 : data <= 8'b00000000 ;
			15'h00004D92 : data <= 8'b00000000 ;
			15'h00004D93 : data <= 8'b00000000 ;
			15'h00004D94 : data <= 8'b00000000 ;
			15'h00004D95 : data <= 8'b00000000 ;
			15'h00004D96 : data <= 8'b00000000 ;
			15'h00004D97 : data <= 8'b00000000 ;
			15'h00004D98 : data <= 8'b00000000 ;
			15'h00004D99 : data <= 8'b00000000 ;
			15'h00004D9A : data <= 8'b00000000 ;
			15'h00004D9B : data <= 8'b00000000 ;
			15'h00004D9C : data <= 8'b00000000 ;
			15'h00004D9D : data <= 8'b00000000 ;
			15'h00004D9E : data <= 8'b00000000 ;
			15'h00004D9F : data <= 8'b00000000 ;
			15'h00004DA0 : data <= 8'b00000000 ;
			15'h00004DA1 : data <= 8'b00000000 ;
			15'h00004DA2 : data <= 8'b00000000 ;
			15'h00004DA3 : data <= 8'b00000000 ;
			15'h00004DA4 : data <= 8'b00000000 ;
			15'h00004DA5 : data <= 8'b00000000 ;
			15'h00004DA6 : data <= 8'b00000000 ;
			15'h00004DA7 : data <= 8'b00000000 ;
			15'h00004DA8 : data <= 8'b00000000 ;
			15'h00004DA9 : data <= 8'b00000000 ;
			15'h00004DAA : data <= 8'b00000000 ;
			15'h00004DAB : data <= 8'b00000000 ;
			15'h00004DAC : data <= 8'b00000000 ;
			15'h00004DAD : data <= 8'b00000000 ;
			15'h00004DAE : data <= 8'b00000000 ;
			15'h00004DAF : data <= 8'b00000000 ;
			15'h00004DB0 : data <= 8'b00000000 ;
			15'h00004DB1 : data <= 8'b00000000 ;
			15'h00004DB2 : data <= 8'b00000000 ;
			15'h00004DB3 : data <= 8'b00000000 ;
			15'h00004DB4 : data <= 8'b00000000 ;
			15'h00004DB5 : data <= 8'b00000000 ;
			15'h00004DB6 : data <= 8'b00000000 ;
			15'h00004DB7 : data <= 8'b00000000 ;
			15'h00004DB8 : data <= 8'b00000000 ;
			15'h00004DB9 : data <= 8'b00000000 ;
			15'h00004DBA : data <= 8'b00000000 ;
			15'h00004DBB : data <= 8'b00000000 ;
			15'h00004DBC : data <= 8'b00000000 ;
			15'h00004DBD : data <= 8'b00000000 ;
			15'h00004DBE : data <= 8'b00000000 ;
			15'h00004DBF : data <= 8'b00000000 ;
			15'h00004DC0 : data <= 8'b00000000 ;
			15'h00004DC1 : data <= 8'b00000000 ;
			15'h00004DC2 : data <= 8'b00000000 ;
			15'h00004DC3 : data <= 8'b00000000 ;
			15'h00004DC4 : data <= 8'b00000000 ;
			15'h00004DC5 : data <= 8'b00000000 ;
			15'h00004DC6 : data <= 8'b00000000 ;
			15'h00004DC7 : data <= 8'b00000000 ;
			15'h00004DC8 : data <= 8'b00000000 ;
			15'h00004DC9 : data <= 8'b00000000 ;
			15'h00004DCA : data <= 8'b00000000 ;
			15'h00004DCB : data <= 8'b00000000 ;
			15'h00004DCC : data <= 8'b00000000 ;
			15'h00004DCD : data <= 8'b00000000 ;
			15'h00004DCE : data <= 8'b00000000 ;
			15'h00004DCF : data <= 8'b00000000 ;
			15'h00004DD0 : data <= 8'b00000000 ;
			15'h00004DD1 : data <= 8'b00000000 ;
			15'h00004DD2 : data <= 8'b00000000 ;
			15'h00004DD3 : data <= 8'b00000000 ;
			15'h00004DD4 : data <= 8'b00000000 ;
			15'h00004DD5 : data <= 8'b00000000 ;
			15'h00004DD6 : data <= 8'b00000000 ;
			15'h00004DD7 : data <= 8'b00000000 ;
			15'h00004DD8 : data <= 8'b00000000 ;
			15'h00004DD9 : data <= 8'b00000000 ;
			15'h00004DDA : data <= 8'b00000000 ;
			15'h00004DDB : data <= 8'b00000000 ;
			15'h00004DDC : data <= 8'b00000000 ;
			15'h00004DDD : data <= 8'b00000000 ;
			15'h00004DDE : data <= 8'b00000000 ;
			15'h00004DDF : data <= 8'b00000000 ;
			15'h00004DE0 : data <= 8'b00000000 ;
			15'h00004DE1 : data <= 8'b00000000 ;
			15'h00004DE2 : data <= 8'b00000000 ;
			15'h00004DE3 : data <= 8'b00000000 ;
			15'h00004DE4 : data <= 8'b00000000 ;
			15'h00004DE5 : data <= 8'b00000000 ;
			15'h00004DE6 : data <= 8'b00000000 ;
			15'h00004DE7 : data <= 8'b00000000 ;
			15'h00004DE8 : data <= 8'b00000000 ;
			15'h00004DE9 : data <= 8'b00000000 ;
			15'h00004DEA : data <= 8'b00000000 ;
			15'h00004DEB : data <= 8'b00000000 ;
			15'h00004DEC : data <= 8'b00000000 ;
			15'h00004DED : data <= 8'b00000000 ;
			15'h00004DEE : data <= 8'b00000000 ;
			15'h00004DEF : data <= 8'b00000000 ;
			15'h00004DF0 : data <= 8'b00000000 ;
			15'h00004DF1 : data <= 8'b00000000 ;
			15'h00004DF2 : data <= 8'b00000000 ;
			15'h00004DF3 : data <= 8'b00000000 ;
			15'h00004DF4 : data <= 8'b00000000 ;
			15'h00004DF5 : data <= 8'b00000000 ;
			15'h00004DF6 : data <= 8'b00000000 ;
			15'h00004DF7 : data <= 8'b00000000 ;
			15'h00004DF8 : data <= 8'b00000000 ;
			15'h00004DF9 : data <= 8'b00000000 ;
			15'h00004DFA : data <= 8'b00000000 ;
			15'h00004DFB : data <= 8'b00000000 ;
			15'h00004DFC : data <= 8'b00000000 ;
			15'h00004DFD : data <= 8'b00000000 ;
			15'h00004DFE : data <= 8'b00000000 ;
			15'h00004DFF : data <= 8'b00000000 ;
			15'h00004E00 : data <= 8'b00000000 ;
			15'h00004E01 : data <= 8'b00000000 ;
			15'h00004E02 : data <= 8'b00000000 ;
			15'h00004E03 : data <= 8'b00000000 ;
			15'h00004E04 : data <= 8'b00000000 ;
			15'h00004E05 : data <= 8'b00000000 ;
			15'h00004E06 : data <= 8'b00000000 ;
			15'h00004E07 : data <= 8'b00000000 ;
			15'h00004E08 : data <= 8'b00000000 ;
			15'h00004E09 : data <= 8'b00000000 ;
			15'h00004E0A : data <= 8'b00000000 ;
			15'h00004E0B : data <= 8'b00000000 ;
			15'h00004E0C : data <= 8'b00000000 ;
			15'h00004E0D : data <= 8'b00000000 ;
			15'h00004E0E : data <= 8'b00000000 ;
			15'h00004E0F : data <= 8'b00000000 ;
			15'h00004E10 : data <= 8'b00000000 ;
			15'h00004E11 : data <= 8'b00000000 ;
			15'h00004E12 : data <= 8'b00000000 ;
			15'h00004E13 : data <= 8'b00000000 ;
			15'h00004E14 : data <= 8'b00000000 ;
			15'h00004E15 : data <= 8'b00000000 ;
			15'h00004E16 : data <= 8'b00000000 ;
			15'h00004E17 : data <= 8'b00000000 ;
			15'h00004E18 : data <= 8'b00000000 ;
			15'h00004E19 : data <= 8'b00000000 ;
			15'h00004E1A : data <= 8'b00000000 ;
			15'h00004E1B : data <= 8'b00000000 ;
			15'h00004E1C : data <= 8'b00000000 ;
			15'h00004E1D : data <= 8'b00000000 ;
			15'h00004E1E : data <= 8'b00000000 ;
			15'h00004E1F : data <= 8'b00000000 ;
			15'h00004E20 : data <= 8'b00000000 ;
			15'h00004E21 : data <= 8'b00000000 ;
			15'h00004E22 : data <= 8'b00000000 ;
			15'h00004E23 : data <= 8'b00000000 ;
			15'h00004E24 : data <= 8'b00000000 ;
			15'h00004E25 : data <= 8'b00000000 ;
			15'h00004E26 : data <= 8'b00000000 ;
			15'h00004E27 : data <= 8'b00000000 ;
			15'h00004E28 : data <= 8'b00000000 ;
			15'h00004E29 : data <= 8'b00000000 ;
			15'h00004E2A : data <= 8'b00000000 ;
			15'h00004E2B : data <= 8'b00000000 ;
			15'h00004E2C : data <= 8'b00000000 ;
			15'h00004E2D : data <= 8'b00000000 ;
			15'h00004E2E : data <= 8'b00000000 ;
			15'h00004E2F : data <= 8'b00000000 ;
			15'h00004E30 : data <= 8'b00000000 ;
			15'h00004E31 : data <= 8'b00000000 ;
			15'h00004E32 : data <= 8'b00000000 ;
			15'h00004E33 : data <= 8'b00000000 ;
			15'h00004E34 : data <= 8'b00000000 ;
			15'h00004E35 : data <= 8'b00000000 ;
			15'h00004E36 : data <= 8'b00000000 ;
			15'h00004E37 : data <= 8'b00000000 ;
			15'h00004E38 : data <= 8'b00000000 ;
			15'h00004E39 : data <= 8'b00000000 ;
			15'h00004E3A : data <= 8'b00000000 ;
			15'h00004E3B : data <= 8'b00000000 ;
			15'h00004E3C : data <= 8'b00000000 ;
			15'h00004E3D : data <= 8'b00000000 ;
			15'h00004E3E : data <= 8'b00000000 ;
			15'h00004E3F : data <= 8'b00000000 ;
			15'h00004E40 : data <= 8'b00000000 ;
			15'h00004E41 : data <= 8'b00000000 ;
			15'h00004E42 : data <= 8'b00000000 ;
			15'h00004E43 : data <= 8'b00000000 ;
			15'h00004E44 : data <= 8'b00000000 ;
			15'h00004E45 : data <= 8'b00000000 ;
			15'h00004E46 : data <= 8'b00000000 ;
			15'h00004E47 : data <= 8'b00000000 ;
			15'h00004E48 : data <= 8'b00000000 ;
			15'h00004E49 : data <= 8'b00000000 ;
			15'h00004E4A : data <= 8'b00000000 ;
			15'h00004E4B : data <= 8'b00000000 ;
			15'h00004E4C : data <= 8'b00000000 ;
			15'h00004E4D : data <= 8'b00000000 ;
			15'h00004E4E : data <= 8'b00000000 ;
			15'h00004E4F : data <= 8'b00000000 ;
			15'h00004E50 : data <= 8'b00000000 ;
			15'h00004E51 : data <= 8'b00000000 ;
			15'h00004E52 : data <= 8'b00000000 ;
			15'h00004E53 : data <= 8'b00000000 ;
			15'h00004E54 : data <= 8'b00000000 ;
			15'h00004E55 : data <= 8'b00000000 ;
			15'h00004E56 : data <= 8'b00000000 ;
			15'h00004E57 : data <= 8'b00000000 ;
			15'h00004E58 : data <= 8'b00000000 ;
			15'h00004E59 : data <= 8'b00000000 ;
			15'h00004E5A : data <= 8'b00000000 ;
			15'h00004E5B : data <= 8'b00000000 ;
			15'h00004E5C : data <= 8'b00000000 ;
			15'h00004E5D : data <= 8'b00000000 ;
			15'h00004E5E : data <= 8'b00000000 ;
			15'h00004E5F : data <= 8'b00000000 ;
			15'h00004E60 : data <= 8'b00000000 ;
			15'h00004E61 : data <= 8'b00000000 ;
			15'h00004E62 : data <= 8'b00000000 ;
			15'h00004E63 : data <= 8'b00000000 ;
			15'h00004E64 : data <= 8'b00000000 ;
			15'h00004E65 : data <= 8'b00000000 ;
			15'h00004E66 : data <= 8'b00000000 ;
			15'h00004E67 : data <= 8'b00000000 ;
			15'h00004E68 : data <= 8'b00000000 ;
			15'h00004E69 : data <= 8'b00000000 ;
			15'h00004E6A : data <= 8'b00000000 ;
			15'h00004E6B : data <= 8'b00000000 ;
			15'h00004E6C : data <= 8'b00000000 ;
			15'h00004E6D : data <= 8'b00000000 ;
			15'h00004E6E : data <= 8'b00000000 ;
			15'h00004E6F : data <= 8'b00000000 ;
			15'h00004E70 : data <= 8'b00000000 ;
			15'h00004E71 : data <= 8'b00000000 ;
			15'h00004E72 : data <= 8'b00000000 ;
			15'h00004E73 : data <= 8'b00000000 ;
			15'h00004E74 : data <= 8'b00000000 ;
			15'h00004E75 : data <= 8'b00000000 ;
			15'h00004E76 : data <= 8'b00000000 ;
			15'h00004E77 : data <= 8'b00000000 ;
			15'h00004E78 : data <= 8'b00000000 ;
			15'h00004E79 : data <= 8'b00000000 ;
			15'h00004E7A : data <= 8'b00000000 ;
			15'h00004E7B : data <= 8'b00000000 ;
			15'h00004E7C : data <= 8'b00000000 ;
			15'h00004E7D : data <= 8'b00000000 ;
			15'h00004E7E : data <= 8'b00000000 ;
			15'h00004E7F : data <= 8'b00000000 ;
			15'h00004E80 : data <= 8'b00000000 ;
			15'h00004E81 : data <= 8'b00000000 ;
			15'h00004E82 : data <= 8'b00000000 ;
			15'h00004E83 : data <= 8'b00000000 ;
			15'h00004E84 : data <= 8'b00000000 ;
			15'h00004E85 : data <= 8'b00000000 ;
			15'h00004E86 : data <= 8'b00000000 ;
			15'h00004E87 : data <= 8'b00000000 ;
			15'h00004E88 : data <= 8'b00000000 ;
			15'h00004E89 : data <= 8'b00000000 ;
			15'h00004E8A : data <= 8'b00000000 ;
			15'h00004E8B : data <= 8'b00000000 ;
			15'h00004E8C : data <= 8'b00000000 ;
			15'h00004E8D : data <= 8'b00000000 ;
			15'h00004E8E : data <= 8'b00000000 ;
			15'h00004E8F : data <= 8'b00000000 ;
			15'h00004E90 : data <= 8'b00000000 ;
			15'h00004E91 : data <= 8'b00000000 ;
			15'h00004E92 : data <= 8'b00000000 ;
			15'h00004E93 : data <= 8'b00000000 ;
			15'h00004E94 : data <= 8'b00000000 ;
			15'h00004E95 : data <= 8'b00000000 ;
			15'h00004E96 : data <= 8'b00000000 ;
			15'h00004E97 : data <= 8'b00000000 ;
			15'h00004E98 : data <= 8'b00000000 ;
			15'h00004E99 : data <= 8'b00000000 ;
			15'h00004E9A : data <= 8'b00000000 ;
			15'h00004E9B : data <= 8'b00000000 ;
			15'h00004E9C : data <= 8'b00000000 ;
			15'h00004E9D : data <= 8'b00000000 ;
			15'h00004E9E : data <= 8'b00000000 ;
			15'h00004E9F : data <= 8'b00000000 ;
			15'h00004EA0 : data <= 8'b00000000 ;
			15'h00004EA1 : data <= 8'b00000000 ;
			15'h00004EA2 : data <= 8'b00000000 ;
			15'h00004EA3 : data <= 8'b00000000 ;
			15'h00004EA4 : data <= 8'b00000000 ;
			15'h00004EA5 : data <= 8'b00000000 ;
			15'h00004EA6 : data <= 8'b00000000 ;
			15'h00004EA7 : data <= 8'b00000000 ;
			15'h00004EA8 : data <= 8'b00000000 ;
			15'h00004EA9 : data <= 8'b00000000 ;
			15'h00004EAA : data <= 8'b00000000 ;
			15'h00004EAB : data <= 8'b00000000 ;
			15'h00004EAC : data <= 8'b00000000 ;
			15'h00004EAD : data <= 8'b00000000 ;
			15'h00004EAE : data <= 8'b00000000 ;
			15'h00004EAF : data <= 8'b00000000 ;
			15'h00004EB0 : data <= 8'b00000000 ;
			15'h00004EB1 : data <= 8'b00000000 ;
			15'h00004EB2 : data <= 8'b00000000 ;
			15'h00004EB3 : data <= 8'b00000000 ;
			15'h00004EB4 : data <= 8'b00000000 ;
			15'h00004EB5 : data <= 8'b00000000 ;
			15'h00004EB6 : data <= 8'b00000000 ;
			15'h00004EB7 : data <= 8'b00000000 ;
			15'h00004EB8 : data <= 8'b00000000 ;
			15'h00004EB9 : data <= 8'b00000000 ;
			15'h00004EBA : data <= 8'b00000000 ;
			15'h00004EBB : data <= 8'b00000000 ;
			15'h00004EBC : data <= 8'b00000000 ;
			15'h00004EBD : data <= 8'b00000000 ;
			15'h00004EBE : data <= 8'b00000000 ;
			15'h00004EBF : data <= 8'b00000000 ;
			15'h00004EC0 : data <= 8'b00000000 ;
			15'h00004EC1 : data <= 8'b00000000 ;
			15'h00004EC2 : data <= 8'b00000000 ;
			15'h00004EC3 : data <= 8'b00000000 ;
			15'h00004EC4 : data <= 8'b00000000 ;
			15'h00004EC5 : data <= 8'b00000000 ;
			15'h00004EC6 : data <= 8'b00000000 ;
			15'h00004EC7 : data <= 8'b00000000 ;
			15'h00004EC8 : data <= 8'b00000000 ;
			15'h00004EC9 : data <= 8'b00000000 ;
			15'h00004ECA : data <= 8'b00000000 ;
			15'h00004ECB : data <= 8'b00000000 ;
			15'h00004ECC : data <= 8'b00000000 ;
			15'h00004ECD : data <= 8'b00000000 ;
			15'h00004ECE : data <= 8'b00000000 ;
			15'h00004ECF : data <= 8'b00000000 ;
			15'h00004ED0 : data <= 8'b00000000 ;
			15'h00004ED1 : data <= 8'b00000000 ;
			15'h00004ED2 : data <= 8'b00000000 ;
			15'h00004ED3 : data <= 8'b00000000 ;
			15'h00004ED4 : data <= 8'b00000000 ;
			15'h00004ED5 : data <= 8'b00000000 ;
			15'h00004ED6 : data <= 8'b00000000 ;
			15'h00004ED7 : data <= 8'b00000000 ;
			15'h00004ED8 : data <= 8'b00000000 ;
			15'h00004ED9 : data <= 8'b00000000 ;
			15'h00004EDA : data <= 8'b00000000 ;
			15'h00004EDB : data <= 8'b00000000 ;
			15'h00004EDC : data <= 8'b00000000 ;
			15'h00004EDD : data <= 8'b00000000 ;
			15'h00004EDE : data <= 8'b00000000 ;
			15'h00004EDF : data <= 8'b00000000 ;
			15'h00004EE0 : data <= 8'b00000000 ;
			15'h00004EE1 : data <= 8'b00000000 ;
			15'h00004EE2 : data <= 8'b00000000 ;
			15'h00004EE3 : data <= 8'b00000000 ;
			15'h00004EE4 : data <= 8'b00000000 ;
			15'h00004EE5 : data <= 8'b00000000 ;
			15'h00004EE6 : data <= 8'b00000000 ;
			15'h00004EE7 : data <= 8'b00000000 ;
			15'h00004EE8 : data <= 8'b00000000 ;
			15'h00004EE9 : data <= 8'b00000000 ;
			15'h00004EEA : data <= 8'b00000000 ;
			15'h00004EEB : data <= 8'b00000000 ;
			15'h00004EEC : data <= 8'b00000000 ;
			15'h00004EED : data <= 8'b00000000 ;
			15'h00004EEE : data <= 8'b00000000 ;
			15'h00004EEF : data <= 8'b00000000 ;
			15'h00004EF0 : data <= 8'b00000000 ;
			15'h00004EF1 : data <= 8'b00000000 ;
			15'h00004EF2 : data <= 8'b00000000 ;
			15'h00004EF3 : data <= 8'b00000000 ;
			15'h00004EF4 : data <= 8'b00000000 ;
			15'h00004EF5 : data <= 8'b00000000 ;
			15'h00004EF6 : data <= 8'b00000000 ;
			15'h00004EF7 : data <= 8'b00000000 ;
			15'h00004EF8 : data <= 8'b00000000 ;
			15'h00004EF9 : data <= 8'b00000000 ;
			15'h00004EFA : data <= 8'b00000000 ;
			15'h00004EFB : data <= 8'b00000000 ;
			15'h00004EFC : data <= 8'b00000000 ;
			15'h00004EFD : data <= 8'b00000000 ;
			15'h00004EFE : data <= 8'b00000000 ;
			15'h00004EFF : data <= 8'b00000000 ;
			15'h00004F00 : data <= 8'b00000000 ;
			15'h00004F01 : data <= 8'b00000000 ;
			15'h00004F02 : data <= 8'b00000000 ;
			15'h00004F03 : data <= 8'b00000000 ;
			15'h00004F04 : data <= 8'b00000000 ;
			15'h00004F05 : data <= 8'b00000000 ;
			15'h00004F06 : data <= 8'b00000000 ;
			15'h00004F07 : data <= 8'b00000000 ;
			15'h00004F08 : data <= 8'b00000000 ;
			15'h00004F09 : data <= 8'b00000000 ;
			15'h00004F0A : data <= 8'b00000000 ;
			15'h00004F0B : data <= 8'b00000000 ;
			15'h00004F0C : data <= 8'b00000000 ;
			15'h00004F0D : data <= 8'b00000000 ;
			15'h00004F0E : data <= 8'b00000000 ;
			15'h00004F0F : data <= 8'b00000000 ;
			15'h00004F10 : data <= 8'b00000000 ;
			15'h00004F11 : data <= 8'b00000000 ;
			15'h00004F12 : data <= 8'b00000000 ;
			15'h00004F13 : data <= 8'b00000000 ;
			15'h00004F14 : data <= 8'b00000000 ;
			15'h00004F15 : data <= 8'b00000000 ;
			15'h00004F16 : data <= 8'b00000000 ;
			15'h00004F17 : data <= 8'b00000000 ;
			15'h00004F18 : data <= 8'b00000000 ;
			15'h00004F19 : data <= 8'b00000000 ;
			15'h00004F1A : data <= 8'b00000000 ;
			15'h00004F1B : data <= 8'b00000000 ;
			15'h00004F1C : data <= 8'b00000000 ;
			15'h00004F1D : data <= 8'b00000000 ;
			15'h00004F1E : data <= 8'b00000000 ;
			15'h00004F1F : data <= 8'b00000000 ;
			15'h00004F20 : data <= 8'b00000000 ;
			15'h00004F21 : data <= 8'b00000000 ;
			15'h00004F22 : data <= 8'b00000000 ;
			15'h00004F23 : data <= 8'b00000000 ;
			15'h00004F24 : data <= 8'b00000000 ;
			15'h00004F25 : data <= 8'b00000000 ;
			15'h00004F26 : data <= 8'b00000000 ;
			15'h00004F27 : data <= 8'b00000000 ;
			15'h00004F28 : data <= 8'b00000000 ;
			15'h00004F29 : data <= 8'b00000000 ;
			15'h00004F2A : data <= 8'b00000000 ;
			15'h00004F2B : data <= 8'b00000000 ;
			15'h00004F2C : data <= 8'b00000000 ;
			15'h00004F2D : data <= 8'b00000000 ;
			15'h00004F2E : data <= 8'b00000000 ;
			15'h00004F2F : data <= 8'b00000000 ;
			15'h00004F30 : data <= 8'b00000000 ;
			15'h00004F31 : data <= 8'b00000000 ;
			15'h00004F32 : data <= 8'b00000000 ;
			15'h00004F33 : data <= 8'b00000000 ;
			15'h00004F34 : data <= 8'b00000000 ;
			15'h00004F35 : data <= 8'b00000000 ;
			15'h00004F36 : data <= 8'b00000000 ;
			15'h00004F37 : data <= 8'b00000000 ;
			15'h00004F38 : data <= 8'b00000000 ;
			15'h00004F39 : data <= 8'b00000000 ;
			15'h00004F3A : data <= 8'b00000000 ;
			15'h00004F3B : data <= 8'b00000000 ;
			15'h00004F3C : data <= 8'b00000000 ;
			15'h00004F3D : data <= 8'b00000000 ;
			15'h00004F3E : data <= 8'b00000000 ;
			15'h00004F3F : data <= 8'b00000000 ;
			15'h00004F40 : data <= 8'b00000000 ;
			15'h00004F41 : data <= 8'b00000000 ;
			15'h00004F42 : data <= 8'b00000000 ;
			15'h00004F43 : data <= 8'b00000000 ;
			15'h00004F44 : data <= 8'b00000000 ;
			15'h00004F45 : data <= 8'b00000000 ;
			15'h00004F46 : data <= 8'b00000000 ;
			15'h00004F47 : data <= 8'b00000000 ;
			15'h00004F48 : data <= 8'b00000000 ;
			15'h00004F49 : data <= 8'b00000000 ;
			15'h00004F4A : data <= 8'b00000000 ;
			15'h00004F4B : data <= 8'b00000000 ;
			15'h00004F4C : data <= 8'b00000000 ;
			15'h00004F4D : data <= 8'b00000000 ;
			15'h00004F4E : data <= 8'b00000000 ;
			15'h00004F4F : data <= 8'b00000000 ;
			15'h00004F50 : data <= 8'b00000000 ;
			15'h00004F51 : data <= 8'b00000000 ;
			15'h00004F52 : data <= 8'b00000000 ;
			15'h00004F53 : data <= 8'b00000000 ;
			15'h00004F54 : data <= 8'b00000000 ;
			15'h00004F55 : data <= 8'b00000000 ;
			15'h00004F56 : data <= 8'b00000000 ;
			15'h00004F57 : data <= 8'b00000000 ;
			15'h00004F58 : data <= 8'b00000000 ;
			15'h00004F59 : data <= 8'b00000000 ;
			15'h00004F5A : data <= 8'b00000000 ;
			15'h00004F5B : data <= 8'b00000000 ;
			15'h00004F5C : data <= 8'b00000000 ;
			15'h00004F5D : data <= 8'b00000000 ;
			15'h00004F5E : data <= 8'b00000000 ;
			15'h00004F5F : data <= 8'b00000000 ;
			15'h00004F60 : data <= 8'b00000000 ;
			15'h00004F61 : data <= 8'b00000000 ;
			15'h00004F62 : data <= 8'b00000000 ;
			15'h00004F63 : data <= 8'b00000000 ;
			15'h00004F64 : data <= 8'b00000000 ;
			15'h00004F65 : data <= 8'b00000000 ;
			15'h00004F66 : data <= 8'b00000000 ;
			15'h00004F67 : data <= 8'b00000000 ;
			15'h00004F68 : data <= 8'b00000000 ;
			15'h00004F69 : data <= 8'b00000000 ;
			15'h00004F6A : data <= 8'b00000000 ;
			15'h00004F6B : data <= 8'b00000000 ;
			15'h00004F6C : data <= 8'b00000000 ;
			15'h00004F6D : data <= 8'b00000000 ;
			15'h00004F6E : data <= 8'b00000000 ;
			15'h00004F6F : data <= 8'b00000000 ;
			15'h00004F70 : data <= 8'b00000000 ;
			15'h00004F71 : data <= 8'b00000000 ;
			15'h00004F72 : data <= 8'b00000000 ;
			15'h00004F73 : data <= 8'b00000000 ;
			15'h00004F74 : data <= 8'b00000000 ;
			15'h00004F75 : data <= 8'b00000000 ;
			15'h00004F76 : data <= 8'b00000000 ;
			15'h00004F77 : data <= 8'b00000000 ;
			15'h00004F78 : data <= 8'b00000000 ;
			15'h00004F79 : data <= 8'b00000000 ;
			15'h00004F7A : data <= 8'b00000000 ;
			15'h00004F7B : data <= 8'b00000000 ;
			15'h00004F7C : data <= 8'b00000000 ;
			15'h00004F7D : data <= 8'b00000000 ;
			15'h00004F7E : data <= 8'b00000000 ;
			15'h00004F7F : data <= 8'b00000000 ;
			15'h00004F80 : data <= 8'b00000000 ;
			15'h00004F81 : data <= 8'b00000000 ;
			15'h00004F82 : data <= 8'b00000000 ;
			15'h00004F83 : data <= 8'b00000000 ;
			15'h00004F84 : data <= 8'b00000000 ;
			15'h00004F85 : data <= 8'b00000000 ;
			15'h00004F86 : data <= 8'b00000000 ;
			15'h00004F87 : data <= 8'b00000000 ;
			15'h00004F88 : data <= 8'b00000000 ;
			15'h00004F89 : data <= 8'b00000000 ;
			15'h00004F8A : data <= 8'b00000000 ;
			15'h00004F8B : data <= 8'b00000000 ;
			15'h00004F8C : data <= 8'b00000000 ;
			15'h00004F8D : data <= 8'b00000000 ;
			15'h00004F8E : data <= 8'b00000000 ;
			15'h00004F8F : data <= 8'b00000000 ;
			15'h00004F90 : data <= 8'b00000000 ;
			15'h00004F91 : data <= 8'b00000000 ;
			15'h00004F92 : data <= 8'b00000000 ;
			15'h00004F93 : data <= 8'b00000000 ;
			15'h00004F94 : data <= 8'b00000000 ;
			15'h00004F95 : data <= 8'b00000000 ;
			15'h00004F96 : data <= 8'b00000000 ;
			15'h00004F97 : data <= 8'b00000000 ;
			15'h00004F98 : data <= 8'b00000000 ;
			15'h00004F99 : data <= 8'b00000000 ;
			15'h00004F9A : data <= 8'b00000000 ;
			15'h00004F9B : data <= 8'b00000000 ;
			15'h00004F9C : data <= 8'b00000000 ;
			15'h00004F9D : data <= 8'b00000000 ;
			15'h00004F9E : data <= 8'b00000000 ;
			15'h00004F9F : data <= 8'b00000000 ;
			15'h00004FA0 : data <= 8'b00000000 ;
			15'h00004FA1 : data <= 8'b00000000 ;
			15'h00004FA2 : data <= 8'b00000000 ;
			15'h00004FA3 : data <= 8'b00000000 ;
			15'h00004FA4 : data <= 8'b00000000 ;
			15'h00004FA5 : data <= 8'b00000000 ;
			15'h00004FA6 : data <= 8'b00000000 ;
			15'h00004FA7 : data <= 8'b00000000 ;
			15'h00004FA8 : data <= 8'b00000000 ;
			15'h00004FA9 : data <= 8'b00000000 ;
			15'h00004FAA : data <= 8'b00000000 ;
			15'h00004FAB : data <= 8'b00000000 ;
			15'h00004FAC : data <= 8'b00000000 ;
			15'h00004FAD : data <= 8'b00000000 ;
			15'h00004FAE : data <= 8'b00000000 ;
			15'h00004FAF : data <= 8'b00000000 ;
			15'h00004FB0 : data <= 8'b00000000 ;
			15'h00004FB1 : data <= 8'b00000000 ;
			15'h00004FB2 : data <= 8'b00000000 ;
			15'h00004FB3 : data <= 8'b00000000 ;
			15'h00004FB4 : data <= 8'b00000000 ;
			15'h00004FB5 : data <= 8'b00000000 ;
			15'h00004FB6 : data <= 8'b00000000 ;
			15'h00004FB7 : data <= 8'b00000000 ;
			15'h00004FB8 : data <= 8'b00000000 ;
			15'h00004FB9 : data <= 8'b00000000 ;
			15'h00004FBA : data <= 8'b00000000 ;
			15'h00004FBB : data <= 8'b00000000 ;
			15'h00004FBC : data <= 8'b00000000 ;
			15'h00004FBD : data <= 8'b00000000 ;
			15'h00004FBE : data <= 8'b00000000 ;
			15'h00004FBF : data <= 8'b00000000 ;
			15'h00004FC0 : data <= 8'b00000000 ;
			15'h00004FC1 : data <= 8'b00000000 ;
			15'h00004FC2 : data <= 8'b00000000 ;
			15'h00004FC3 : data <= 8'b00000000 ;
			15'h00004FC4 : data <= 8'b00000000 ;
			15'h00004FC5 : data <= 8'b00000000 ;
			15'h00004FC6 : data <= 8'b00000000 ;
			15'h00004FC7 : data <= 8'b00000000 ;
			15'h00004FC8 : data <= 8'b00000000 ;
			15'h00004FC9 : data <= 8'b00000000 ;
			15'h00004FCA : data <= 8'b00000000 ;
			15'h00004FCB : data <= 8'b00000000 ;
			15'h00004FCC : data <= 8'b00000000 ;
			15'h00004FCD : data <= 8'b00000000 ;
			15'h00004FCE : data <= 8'b00000000 ;
			15'h00004FCF : data <= 8'b00000000 ;
			15'h00004FD0 : data <= 8'b00000000 ;
			15'h00004FD1 : data <= 8'b00000000 ;
			15'h00004FD2 : data <= 8'b00000000 ;
			15'h00004FD3 : data <= 8'b00000000 ;
			15'h00004FD4 : data <= 8'b00000000 ;
			15'h00004FD5 : data <= 8'b00000000 ;
			15'h00004FD6 : data <= 8'b00000000 ;
			15'h00004FD7 : data <= 8'b00000000 ;
			15'h00004FD8 : data <= 8'b00000000 ;
			15'h00004FD9 : data <= 8'b00000000 ;
			15'h00004FDA : data <= 8'b00000000 ;
			15'h00004FDB : data <= 8'b00000000 ;
			15'h00004FDC : data <= 8'b00000000 ;
			15'h00004FDD : data <= 8'b00000000 ;
			15'h00004FDE : data <= 8'b00000000 ;
			15'h00004FDF : data <= 8'b00000000 ;
			15'h00004FE0 : data <= 8'b00000000 ;
			15'h00004FE1 : data <= 8'b00000000 ;
			15'h00004FE2 : data <= 8'b00000000 ;
			15'h00004FE3 : data <= 8'b00000000 ;
			15'h00004FE4 : data <= 8'b00000000 ;
			15'h00004FE5 : data <= 8'b00000000 ;
			15'h00004FE6 : data <= 8'b00000000 ;
			15'h00004FE7 : data <= 8'b00000000 ;
			15'h00004FE8 : data <= 8'b00000000 ;
			15'h00004FE9 : data <= 8'b00000000 ;
			15'h00004FEA : data <= 8'b00000000 ;
			15'h00004FEB : data <= 8'b00000000 ;
			15'h00004FEC : data <= 8'b00000000 ;
			15'h00004FED : data <= 8'b00000000 ;
			15'h00004FEE : data <= 8'b00000000 ;
			15'h00004FEF : data <= 8'b00000000 ;
			15'h00004FF0 : data <= 8'b00000000 ;
			15'h00004FF1 : data <= 8'b00000000 ;
			15'h00004FF2 : data <= 8'b00000000 ;
			15'h00004FF3 : data <= 8'b00000000 ;
			15'h00004FF4 : data <= 8'b00000000 ;
			15'h00004FF5 : data <= 8'b00000000 ;
			15'h00004FF6 : data <= 8'b00000000 ;
			15'h00004FF7 : data <= 8'b00000000 ;
			15'h00004FF8 : data <= 8'b00000000 ;
			15'h00004FF9 : data <= 8'b00000000 ;
			15'h00004FFA : data <= 8'b00000000 ;
			15'h00004FFB : data <= 8'b00000000 ;
			15'h00004FFC : data <= 8'b00000000 ;
			15'h00004FFD : data <= 8'b00000000 ;
			15'h00004FFE : data <= 8'b00000000 ;
			15'h00004FFF : data <= 8'b00000000 ;
			15'h00005000 : data <= 8'b00000000 ;
			15'h00005001 : data <= 8'b00000000 ;
			15'h00005002 : data <= 8'b00000000 ;
			15'h00005003 : data <= 8'b00000000 ;
			15'h00005004 : data <= 8'b00000000 ;
			15'h00005005 : data <= 8'b00000000 ;
			15'h00005006 : data <= 8'b00000000 ;
			15'h00005007 : data <= 8'b00000000 ;
			15'h00005008 : data <= 8'b00000000 ;
			15'h00005009 : data <= 8'b00000000 ;
			15'h0000500A : data <= 8'b00000000 ;
			15'h0000500B : data <= 8'b00000000 ;
			15'h0000500C : data <= 8'b00000000 ;
			15'h0000500D : data <= 8'b00000000 ;
			15'h0000500E : data <= 8'b00000000 ;
			15'h0000500F : data <= 8'b00000000 ;
			15'h00005010 : data <= 8'b00000000 ;
			15'h00005011 : data <= 8'b00000000 ;
			15'h00005012 : data <= 8'b00000000 ;
			15'h00005013 : data <= 8'b00000000 ;
			15'h00005014 : data <= 8'b00000000 ;
			15'h00005015 : data <= 8'b00000000 ;
			15'h00005016 : data <= 8'b00000000 ;
			15'h00005017 : data <= 8'b00000000 ;
			15'h00005018 : data <= 8'b00000000 ;
			15'h00005019 : data <= 8'b00000000 ;
			15'h0000501A : data <= 8'b00000000 ;
			15'h0000501B : data <= 8'b00000000 ;
			15'h0000501C : data <= 8'b00000000 ;
			15'h0000501D : data <= 8'b00000000 ;
			15'h0000501E : data <= 8'b00000000 ;
			15'h0000501F : data <= 8'b00000000 ;
			15'h00005020 : data <= 8'b00000000 ;
			15'h00005021 : data <= 8'b00000000 ;
			15'h00005022 : data <= 8'b00000000 ;
			15'h00005023 : data <= 8'b00000000 ;
			15'h00005024 : data <= 8'b00000000 ;
			15'h00005025 : data <= 8'b00000000 ;
			15'h00005026 : data <= 8'b00000000 ;
			15'h00005027 : data <= 8'b00000000 ;
			15'h00005028 : data <= 8'b00000000 ;
			15'h00005029 : data <= 8'b00000000 ;
			15'h0000502A : data <= 8'b00000000 ;
			15'h0000502B : data <= 8'b00000000 ;
			15'h0000502C : data <= 8'b00000000 ;
			15'h0000502D : data <= 8'b00000000 ;
			15'h0000502E : data <= 8'b00000000 ;
			15'h0000502F : data <= 8'b00000000 ;
			15'h00005030 : data <= 8'b00000000 ;
			15'h00005031 : data <= 8'b00000000 ;
			15'h00005032 : data <= 8'b00000000 ;
			15'h00005033 : data <= 8'b00000000 ;
			15'h00005034 : data <= 8'b00000000 ;
			15'h00005035 : data <= 8'b00000000 ;
			15'h00005036 : data <= 8'b00000000 ;
			15'h00005037 : data <= 8'b00000000 ;
			15'h00005038 : data <= 8'b00000000 ;
			15'h00005039 : data <= 8'b00000000 ;
			15'h0000503A : data <= 8'b00000000 ;
			15'h0000503B : data <= 8'b00000000 ;
			15'h0000503C : data <= 8'b00000000 ;
			15'h0000503D : data <= 8'b00000000 ;
			15'h0000503E : data <= 8'b00000000 ;
			15'h0000503F : data <= 8'b00000000 ;
			15'h00005040 : data <= 8'b00000000 ;
			15'h00005041 : data <= 8'b00000000 ;
			15'h00005042 : data <= 8'b00000000 ;
			15'h00005043 : data <= 8'b00000000 ;
			15'h00005044 : data <= 8'b00000000 ;
			15'h00005045 : data <= 8'b00000000 ;
			15'h00005046 : data <= 8'b00000000 ;
			15'h00005047 : data <= 8'b00000000 ;
			15'h00005048 : data <= 8'b00000000 ;
			15'h00005049 : data <= 8'b00000000 ;
			15'h0000504A : data <= 8'b00000000 ;
			15'h0000504B : data <= 8'b00000000 ;
			15'h0000504C : data <= 8'b00000000 ;
			15'h0000504D : data <= 8'b00000000 ;
			15'h0000504E : data <= 8'b00000000 ;
			15'h0000504F : data <= 8'b00000000 ;
			15'h00005050 : data <= 8'b00000000 ;
			15'h00005051 : data <= 8'b00000000 ;
			15'h00005052 : data <= 8'b00000000 ;
			15'h00005053 : data <= 8'b00000000 ;
			15'h00005054 : data <= 8'b00000000 ;
			15'h00005055 : data <= 8'b00000000 ;
			15'h00005056 : data <= 8'b00000000 ;
			15'h00005057 : data <= 8'b00000000 ;
			15'h00005058 : data <= 8'b00000000 ;
			15'h00005059 : data <= 8'b00000000 ;
			15'h0000505A : data <= 8'b00000000 ;
			15'h0000505B : data <= 8'b00000000 ;
			15'h0000505C : data <= 8'b00000000 ;
			15'h0000505D : data <= 8'b00000000 ;
			15'h0000505E : data <= 8'b00000000 ;
			15'h0000505F : data <= 8'b00000000 ;
			15'h00005060 : data <= 8'b00000000 ;
			15'h00005061 : data <= 8'b00000000 ;
			15'h00005062 : data <= 8'b00000000 ;
			15'h00005063 : data <= 8'b00000000 ;
			15'h00005064 : data <= 8'b00000000 ;
			15'h00005065 : data <= 8'b00000000 ;
			15'h00005066 : data <= 8'b00000000 ;
			15'h00005067 : data <= 8'b00000000 ;
			15'h00005068 : data <= 8'b00000000 ;
			15'h00005069 : data <= 8'b00000000 ;
			15'h0000506A : data <= 8'b00000000 ;
			15'h0000506B : data <= 8'b00000000 ;
			15'h0000506C : data <= 8'b00000000 ;
			15'h0000506D : data <= 8'b00000000 ;
			15'h0000506E : data <= 8'b00000000 ;
			15'h0000506F : data <= 8'b00000000 ;
			15'h00005070 : data <= 8'b00000000 ;
			15'h00005071 : data <= 8'b00000000 ;
			15'h00005072 : data <= 8'b00000000 ;
			15'h00005073 : data <= 8'b00000000 ;
			15'h00005074 : data <= 8'b00000000 ;
			15'h00005075 : data <= 8'b00000000 ;
			15'h00005076 : data <= 8'b00000000 ;
			15'h00005077 : data <= 8'b00000000 ;
			15'h00005078 : data <= 8'b00000000 ;
			15'h00005079 : data <= 8'b00000000 ;
			15'h0000507A : data <= 8'b00000000 ;
			15'h0000507B : data <= 8'b00000000 ;
			15'h0000507C : data <= 8'b00000000 ;
			15'h0000507D : data <= 8'b00000000 ;
			15'h0000507E : data <= 8'b00000000 ;
			15'h0000507F : data <= 8'b00000000 ;
			15'h00005080 : data <= 8'b00000000 ;
			15'h00005081 : data <= 8'b00000000 ;
			15'h00005082 : data <= 8'b00000000 ;
			15'h00005083 : data <= 8'b00000000 ;
			15'h00005084 : data <= 8'b00000000 ;
			15'h00005085 : data <= 8'b00000000 ;
			15'h00005086 : data <= 8'b00000000 ;
			15'h00005087 : data <= 8'b00000000 ;
			15'h00005088 : data <= 8'b00000000 ;
			15'h00005089 : data <= 8'b00000000 ;
			15'h0000508A : data <= 8'b00000000 ;
			15'h0000508B : data <= 8'b00000000 ;
			15'h0000508C : data <= 8'b00000000 ;
			15'h0000508D : data <= 8'b00000000 ;
			15'h0000508E : data <= 8'b00000000 ;
			15'h0000508F : data <= 8'b00000000 ;
			15'h00005090 : data <= 8'b00000000 ;
			15'h00005091 : data <= 8'b00000000 ;
			15'h00005092 : data <= 8'b00000000 ;
			15'h00005093 : data <= 8'b00000000 ;
			15'h00005094 : data <= 8'b00000000 ;
			15'h00005095 : data <= 8'b00000000 ;
			15'h00005096 : data <= 8'b00000000 ;
			15'h00005097 : data <= 8'b00000000 ;
			15'h00005098 : data <= 8'b00000000 ;
			15'h00005099 : data <= 8'b00000000 ;
			15'h0000509A : data <= 8'b00000000 ;
			15'h0000509B : data <= 8'b00000000 ;
			15'h0000509C : data <= 8'b00000000 ;
			15'h0000509D : data <= 8'b00000000 ;
			15'h0000509E : data <= 8'b00000000 ;
			15'h0000509F : data <= 8'b00000000 ;
			15'h000050A0 : data <= 8'b00000000 ;
			15'h000050A1 : data <= 8'b00000000 ;
			15'h000050A2 : data <= 8'b00000000 ;
			15'h000050A3 : data <= 8'b00000000 ;
			15'h000050A4 : data <= 8'b00000000 ;
			15'h000050A5 : data <= 8'b00000000 ;
			15'h000050A6 : data <= 8'b00000000 ;
			15'h000050A7 : data <= 8'b00000000 ;
			15'h000050A8 : data <= 8'b00000000 ;
			15'h000050A9 : data <= 8'b00000000 ;
			15'h000050AA : data <= 8'b00000000 ;
			15'h000050AB : data <= 8'b00000000 ;
			15'h000050AC : data <= 8'b00000000 ;
			15'h000050AD : data <= 8'b00000000 ;
			15'h000050AE : data <= 8'b00000000 ;
			15'h000050AF : data <= 8'b00000000 ;
			15'h000050B0 : data <= 8'b00000000 ;
			15'h000050B1 : data <= 8'b00000000 ;
			15'h000050B2 : data <= 8'b00000000 ;
			15'h000050B3 : data <= 8'b00000000 ;
			15'h000050B4 : data <= 8'b00000000 ;
			15'h000050B5 : data <= 8'b00000000 ;
			15'h000050B6 : data <= 8'b00000000 ;
			15'h000050B7 : data <= 8'b00000000 ;
			15'h000050B8 : data <= 8'b00000000 ;
			15'h000050B9 : data <= 8'b00000000 ;
			15'h000050BA : data <= 8'b00000000 ;
			15'h000050BB : data <= 8'b00000000 ;
			15'h000050BC : data <= 8'b00000000 ;
			15'h000050BD : data <= 8'b00000000 ;
			15'h000050BE : data <= 8'b00000000 ;
			15'h000050BF : data <= 8'b00000000 ;
			15'h000050C0 : data <= 8'b00000000 ;
			15'h000050C1 : data <= 8'b00000000 ;
			15'h000050C2 : data <= 8'b00000000 ;
			15'h000050C3 : data <= 8'b00000000 ;
			15'h000050C4 : data <= 8'b00000000 ;
			15'h000050C5 : data <= 8'b00000000 ;
			15'h000050C6 : data <= 8'b00000000 ;
			15'h000050C7 : data <= 8'b00000000 ;
			15'h000050C8 : data <= 8'b00000000 ;
			15'h000050C9 : data <= 8'b00000000 ;
			15'h000050CA : data <= 8'b00000000 ;
			15'h000050CB : data <= 8'b00000000 ;
			15'h000050CC : data <= 8'b00000000 ;
			15'h000050CD : data <= 8'b00000000 ;
			15'h000050CE : data <= 8'b00000000 ;
			15'h000050CF : data <= 8'b00000000 ;
			15'h000050D0 : data <= 8'b00000000 ;
			15'h000050D1 : data <= 8'b00000000 ;
			15'h000050D2 : data <= 8'b00000000 ;
			15'h000050D3 : data <= 8'b00000000 ;
			15'h000050D4 : data <= 8'b00000000 ;
			15'h000050D5 : data <= 8'b00000000 ;
			15'h000050D6 : data <= 8'b00000000 ;
			15'h000050D7 : data <= 8'b00000000 ;
			15'h000050D8 : data <= 8'b00000000 ;
			15'h000050D9 : data <= 8'b00000000 ;
			15'h000050DA : data <= 8'b00000000 ;
			15'h000050DB : data <= 8'b00000000 ;
			15'h000050DC : data <= 8'b00000000 ;
			15'h000050DD : data <= 8'b00000000 ;
			15'h000050DE : data <= 8'b00000000 ;
			15'h000050DF : data <= 8'b00000000 ;
			15'h000050E0 : data <= 8'b00000000 ;
			15'h000050E1 : data <= 8'b00000000 ;
			15'h000050E2 : data <= 8'b00000000 ;
			15'h000050E3 : data <= 8'b00000000 ;
			15'h000050E4 : data <= 8'b00000000 ;
			15'h000050E5 : data <= 8'b00000000 ;
			15'h000050E6 : data <= 8'b00000000 ;
			15'h000050E7 : data <= 8'b00000000 ;
			15'h000050E8 : data <= 8'b00000000 ;
			15'h000050E9 : data <= 8'b00000000 ;
			15'h000050EA : data <= 8'b00000000 ;
			15'h000050EB : data <= 8'b00000000 ;
			15'h000050EC : data <= 8'b00000000 ;
			15'h000050ED : data <= 8'b00000000 ;
			15'h000050EE : data <= 8'b00000000 ;
			15'h000050EF : data <= 8'b00000000 ;
			15'h000050F0 : data <= 8'b00000000 ;
			15'h000050F1 : data <= 8'b00000000 ;
			15'h000050F2 : data <= 8'b00000000 ;
			15'h000050F3 : data <= 8'b00000000 ;
			15'h000050F4 : data <= 8'b00000000 ;
			15'h000050F5 : data <= 8'b00000000 ;
			15'h000050F6 : data <= 8'b00000000 ;
			15'h000050F7 : data <= 8'b00000000 ;
			15'h000050F8 : data <= 8'b00000000 ;
			15'h000050F9 : data <= 8'b00000000 ;
			15'h000050FA : data <= 8'b00000000 ;
			15'h000050FB : data <= 8'b00000000 ;
			15'h000050FC : data <= 8'b00000000 ;
			15'h000050FD : data <= 8'b00000000 ;
			15'h000050FE : data <= 8'b00000000 ;
			15'h000050FF : data <= 8'b00000000 ;
			15'h00005100 : data <= 8'b00000000 ;
			15'h00005101 : data <= 8'b00000000 ;
			15'h00005102 : data <= 8'b00000000 ;
			15'h00005103 : data <= 8'b00000000 ;
			15'h00005104 : data <= 8'b00000000 ;
			15'h00005105 : data <= 8'b00000000 ;
			15'h00005106 : data <= 8'b00000000 ;
			15'h00005107 : data <= 8'b00000000 ;
			15'h00005108 : data <= 8'b00000000 ;
			15'h00005109 : data <= 8'b00000000 ;
			15'h0000510A : data <= 8'b00000000 ;
			15'h0000510B : data <= 8'b00000000 ;
			15'h0000510C : data <= 8'b00000000 ;
			15'h0000510D : data <= 8'b00000000 ;
			15'h0000510E : data <= 8'b00000000 ;
			15'h0000510F : data <= 8'b00000000 ;
			15'h00005110 : data <= 8'b00000000 ;
			15'h00005111 : data <= 8'b00000000 ;
			15'h00005112 : data <= 8'b00000000 ;
			15'h00005113 : data <= 8'b00000000 ;
			15'h00005114 : data <= 8'b00000000 ;
			15'h00005115 : data <= 8'b00000000 ;
			15'h00005116 : data <= 8'b00000000 ;
			15'h00005117 : data <= 8'b00000000 ;
			15'h00005118 : data <= 8'b00000000 ;
			15'h00005119 : data <= 8'b00000000 ;
			15'h0000511A : data <= 8'b00000000 ;
			15'h0000511B : data <= 8'b00000000 ;
			15'h0000511C : data <= 8'b00000000 ;
			15'h0000511D : data <= 8'b00000000 ;
			15'h0000511E : data <= 8'b00000000 ;
			15'h0000511F : data <= 8'b00000000 ;
			15'h00005120 : data <= 8'b00000000 ;
			15'h00005121 : data <= 8'b00000000 ;
			15'h00005122 : data <= 8'b00000000 ;
			15'h00005123 : data <= 8'b00000000 ;
			15'h00005124 : data <= 8'b00000000 ;
			15'h00005125 : data <= 8'b00000000 ;
			15'h00005126 : data <= 8'b00000000 ;
			15'h00005127 : data <= 8'b00000000 ;
			15'h00005128 : data <= 8'b00000000 ;
			15'h00005129 : data <= 8'b00000000 ;
			15'h0000512A : data <= 8'b00000000 ;
			15'h0000512B : data <= 8'b00000000 ;
			15'h0000512C : data <= 8'b00000000 ;
			15'h0000512D : data <= 8'b00000000 ;
			15'h0000512E : data <= 8'b00000000 ;
			15'h0000512F : data <= 8'b00000000 ;
			15'h00005130 : data <= 8'b00000000 ;
			15'h00005131 : data <= 8'b00000000 ;
			15'h00005132 : data <= 8'b00000000 ;
			15'h00005133 : data <= 8'b00000000 ;
			15'h00005134 : data <= 8'b00000000 ;
			15'h00005135 : data <= 8'b00000000 ;
			15'h00005136 : data <= 8'b00000000 ;
			15'h00005137 : data <= 8'b00000000 ;
			15'h00005138 : data <= 8'b00000000 ;
			15'h00005139 : data <= 8'b00000000 ;
			15'h0000513A : data <= 8'b00000000 ;
			15'h0000513B : data <= 8'b00000000 ;
			15'h0000513C : data <= 8'b00000000 ;
			15'h0000513D : data <= 8'b00000000 ;
			15'h0000513E : data <= 8'b00000000 ;
			15'h0000513F : data <= 8'b00000000 ;
			15'h00005140 : data <= 8'b00000000 ;
			15'h00005141 : data <= 8'b00000000 ;
			15'h00005142 : data <= 8'b00000000 ;
			15'h00005143 : data <= 8'b00000000 ;
			15'h00005144 : data <= 8'b00000000 ;
			15'h00005145 : data <= 8'b00000000 ;
			15'h00005146 : data <= 8'b00000000 ;
			15'h00005147 : data <= 8'b00000000 ;
			15'h00005148 : data <= 8'b00000000 ;
			15'h00005149 : data <= 8'b00000000 ;
			15'h0000514A : data <= 8'b00000000 ;
			15'h0000514B : data <= 8'b00000000 ;
			15'h0000514C : data <= 8'b00000000 ;
			15'h0000514D : data <= 8'b00000000 ;
			15'h0000514E : data <= 8'b00000000 ;
			15'h0000514F : data <= 8'b00000000 ;
			15'h00005150 : data <= 8'b00000000 ;
			15'h00005151 : data <= 8'b00000000 ;
			15'h00005152 : data <= 8'b00000000 ;
			15'h00005153 : data <= 8'b00000000 ;
			15'h00005154 : data <= 8'b00000000 ;
			15'h00005155 : data <= 8'b00000000 ;
			15'h00005156 : data <= 8'b00000000 ;
			15'h00005157 : data <= 8'b00000000 ;
			15'h00005158 : data <= 8'b00000000 ;
			15'h00005159 : data <= 8'b00000000 ;
			15'h0000515A : data <= 8'b00000000 ;
			15'h0000515B : data <= 8'b00000000 ;
			15'h0000515C : data <= 8'b00000000 ;
			15'h0000515D : data <= 8'b00000000 ;
			15'h0000515E : data <= 8'b00000000 ;
			15'h0000515F : data <= 8'b00000000 ;
			15'h00005160 : data <= 8'b00000000 ;
			15'h00005161 : data <= 8'b00000000 ;
			15'h00005162 : data <= 8'b00000000 ;
			15'h00005163 : data <= 8'b00000000 ;
			15'h00005164 : data <= 8'b00000000 ;
			15'h00005165 : data <= 8'b00000000 ;
			15'h00005166 : data <= 8'b00000000 ;
			15'h00005167 : data <= 8'b00000000 ;
			15'h00005168 : data <= 8'b00000000 ;
			15'h00005169 : data <= 8'b00000000 ;
			15'h0000516A : data <= 8'b00000000 ;
			15'h0000516B : data <= 8'b00000000 ;
			15'h0000516C : data <= 8'b00000000 ;
			15'h0000516D : data <= 8'b00000000 ;
			15'h0000516E : data <= 8'b00000000 ;
			15'h0000516F : data <= 8'b00000000 ;
			15'h00005170 : data <= 8'b00000000 ;
			15'h00005171 : data <= 8'b00000000 ;
			15'h00005172 : data <= 8'b00000000 ;
			15'h00005173 : data <= 8'b00000000 ;
			15'h00005174 : data <= 8'b00000000 ;
			15'h00005175 : data <= 8'b00000000 ;
			15'h00005176 : data <= 8'b00000000 ;
			15'h00005177 : data <= 8'b00000000 ;
			15'h00005178 : data <= 8'b00000000 ;
			15'h00005179 : data <= 8'b00000000 ;
			15'h0000517A : data <= 8'b00000000 ;
			15'h0000517B : data <= 8'b00000000 ;
			15'h0000517C : data <= 8'b00000000 ;
			15'h0000517D : data <= 8'b00000000 ;
			15'h0000517E : data <= 8'b00000000 ;
			15'h0000517F : data <= 8'b00000000 ;
			15'h00005180 : data <= 8'b00000000 ;
			15'h00005181 : data <= 8'b00000000 ;
			15'h00005182 : data <= 8'b00000000 ;
			15'h00005183 : data <= 8'b00000000 ;
			15'h00005184 : data <= 8'b00000000 ;
			15'h00005185 : data <= 8'b00000000 ;
			15'h00005186 : data <= 8'b00000000 ;
			15'h00005187 : data <= 8'b00000000 ;
			15'h00005188 : data <= 8'b00000000 ;
			15'h00005189 : data <= 8'b00000000 ;
			15'h0000518A : data <= 8'b00000000 ;
			15'h0000518B : data <= 8'b00000000 ;
			15'h0000518C : data <= 8'b00000000 ;
			15'h0000518D : data <= 8'b00000000 ;
			15'h0000518E : data <= 8'b00000000 ;
			15'h0000518F : data <= 8'b00000000 ;
			15'h00005190 : data <= 8'b00000000 ;
			15'h00005191 : data <= 8'b00000000 ;
			15'h00005192 : data <= 8'b00000000 ;
			15'h00005193 : data <= 8'b00000000 ;
			15'h00005194 : data <= 8'b00000000 ;
			15'h00005195 : data <= 8'b00000000 ;
			15'h00005196 : data <= 8'b00000000 ;
			15'h00005197 : data <= 8'b00000000 ;
			15'h00005198 : data <= 8'b00000000 ;
			15'h00005199 : data <= 8'b00000000 ;
			15'h0000519A : data <= 8'b00000000 ;
			15'h0000519B : data <= 8'b00000000 ;
			15'h0000519C : data <= 8'b00000000 ;
			15'h0000519D : data <= 8'b00000000 ;
			15'h0000519E : data <= 8'b00000000 ;
			15'h0000519F : data <= 8'b00000000 ;
			15'h000051A0 : data <= 8'b00000000 ;
			15'h000051A1 : data <= 8'b00000000 ;
			15'h000051A2 : data <= 8'b00000000 ;
			15'h000051A3 : data <= 8'b00000000 ;
			15'h000051A4 : data <= 8'b00000000 ;
			15'h000051A5 : data <= 8'b00000000 ;
			15'h000051A6 : data <= 8'b00000000 ;
			15'h000051A7 : data <= 8'b00000000 ;
			15'h000051A8 : data <= 8'b00000000 ;
			15'h000051A9 : data <= 8'b00000000 ;
			15'h000051AA : data <= 8'b00000000 ;
			15'h000051AB : data <= 8'b00000000 ;
			15'h000051AC : data <= 8'b00000000 ;
			15'h000051AD : data <= 8'b00000000 ;
			15'h000051AE : data <= 8'b00000000 ;
			15'h000051AF : data <= 8'b00000000 ;
			15'h000051B0 : data <= 8'b00000000 ;
			15'h000051B1 : data <= 8'b00000000 ;
			15'h000051B2 : data <= 8'b00000000 ;
			15'h000051B3 : data <= 8'b00000000 ;
			15'h000051B4 : data <= 8'b00000000 ;
			15'h000051B5 : data <= 8'b00000000 ;
			15'h000051B6 : data <= 8'b00000000 ;
			15'h000051B7 : data <= 8'b00000000 ;
			15'h000051B8 : data <= 8'b00000000 ;
			15'h000051B9 : data <= 8'b00000000 ;
			15'h000051BA : data <= 8'b00000000 ;
			15'h000051BB : data <= 8'b00000000 ;
			15'h000051BC : data <= 8'b00000000 ;
			15'h000051BD : data <= 8'b00000000 ;
			15'h000051BE : data <= 8'b00000000 ;
			15'h000051BF : data <= 8'b00000000 ;
			15'h000051C0 : data <= 8'b00000000 ;
			15'h000051C1 : data <= 8'b00000000 ;
			15'h000051C2 : data <= 8'b00000000 ;
			15'h000051C3 : data <= 8'b00000000 ;
			15'h000051C4 : data <= 8'b00000000 ;
			15'h000051C5 : data <= 8'b00000000 ;
			15'h000051C6 : data <= 8'b00000000 ;
			15'h000051C7 : data <= 8'b00000000 ;
			15'h000051C8 : data <= 8'b00000000 ;
			15'h000051C9 : data <= 8'b00000000 ;
			15'h000051CA : data <= 8'b00000000 ;
			15'h000051CB : data <= 8'b00000000 ;
			15'h000051CC : data <= 8'b00000000 ;
			15'h000051CD : data <= 8'b00000000 ;
			15'h000051CE : data <= 8'b00000000 ;
			15'h000051CF : data <= 8'b00000000 ;
			15'h000051D0 : data <= 8'b00000000 ;
			15'h000051D1 : data <= 8'b00000000 ;
			15'h000051D2 : data <= 8'b00000000 ;
			15'h000051D3 : data <= 8'b00000000 ;
			15'h000051D4 : data <= 8'b00000000 ;
			15'h000051D5 : data <= 8'b00000000 ;
			15'h000051D6 : data <= 8'b00000000 ;
			15'h000051D7 : data <= 8'b00000000 ;
			15'h000051D8 : data <= 8'b00000000 ;
			15'h000051D9 : data <= 8'b00000000 ;
			15'h000051DA : data <= 8'b00000000 ;
			15'h000051DB : data <= 8'b00000000 ;
			15'h000051DC : data <= 8'b00000000 ;
			15'h000051DD : data <= 8'b00000000 ;
			15'h000051DE : data <= 8'b00000000 ;
			15'h000051DF : data <= 8'b00000000 ;
			15'h000051E0 : data <= 8'b00000000 ;
			15'h000051E1 : data <= 8'b00000000 ;
			15'h000051E2 : data <= 8'b00000000 ;
			15'h000051E3 : data <= 8'b00000000 ;
			15'h000051E4 : data <= 8'b00000000 ;
			15'h000051E5 : data <= 8'b00000000 ;
			15'h000051E6 : data <= 8'b00000000 ;
			15'h000051E7 : data <= 8'b00000000 ;
			15'h000051E8 : data <= 8'b00000000 ;
			15'h000051E9 : data <= 8'b00000000 ;
			15'h000051EA : data <= 8'b00000000 ;
			15'h000051EB : data <= 8'b00000000 ;
			15'h000051EC : data <= 8'b00000000 ;
			15'h000051ED : data <= 8'b00000000 ;
			15'h000051EE : data <= 8'b00000000 ;
			15'h000051EF : data <= 8'b00000000 ;
			15'h000051F0 : data <= 8'b00000000 ;
			15'h000051F1 : data <= 8'b00000000 ;
			15'h000051F2 : data <= 8'b00000000 ;
			15'h000051F3 : data <= 8'b00000000 ;
			15'h000051F4 : data <= 8'b00000000 ;
			15'h000051F5 : data <= 8'b00000000 ;
			15'h000051F6 : data <= 8'b00000000 ;
			15'h000051F7 : data <= 8'b00000000 ;
			15'h000051F8 : data <= 8'b00000000 ;
			15'h000051F9 : data <= 8'b00000000 ;
			15'h000051FA : data <= 8'b00000000 ;
			15'h000051FB : data <= 8'b00000000 ;
			15'h000051FC : data <= 8'b00000000 ;
			15'h000051FD : data <= 8'b00000000 ;
			15'h000051FE : data <= 8'b00000000 ;
			15'h000051FF : data <= 8'b00000000 ;
			15'h00005200 : data <= 8'b00000000 ;
			15'h00005201 : data <= 8'b00000000 ;
			15'h00005202 : data <= 8'b00000000 ;
			15'h00005203 : data <= 8'b00000000 ;
			15'h00005204 : data <= 8'b00000000 ;
			15'h00005205 : data <= 8'b00000000 ;
			15'h00005206 : data <= 8'b00000000 ;
			15'h00005207 : data <= 8'b00000000 ;
			15'h00005208 : data <= 8'b00000000 ;
			15'h00005209 : data <= 8'b00000000 ;
			15'h0000520A : data <= 8'b00000000 ;
			15'h0000520B : data <= 8'b00000000 ;
			15'h0000520C : data <= 8'b00000000 ;
			15'h0000520D : data <= 8'b00000000 ;
			15'h0000520E : data <= 8'b00000000 ;
			15'h0000520F : data <= 8'b00000000 ;
			15'h00005210 : data <= 8'b00000000 ;
			15'h00005211 : data <= 8'b00000000 ;
			15'h00005212 : data <= 8'b00000000 ;
			15'h00005213 : data <= 8'b00000000 ;
			15'h00005214 : data <= 8'b00000000 ;
			15'h00005215 : data <= 8'b00000000 ;
			15'h00005216 : data <= 8'b00000000 ;
			15'h00005217 : data <= 8'b00000000 ;
			15'h00005218 : data <= 8'b00000000 ;
			15'h00005219 : data <= 8'b00000000 ;
			15'h0000521A : data <= 8'b00000000 ;
			15'h0000521B : data <= 8'b00000000 ;
			15'h0000521C : data <= 8'b00000000 ;
			15'h0000521D : data <= 8'b00000000 ;
			15'h0000521E : data <= 8'b00000000 ;
			15'h0000521F : data <= 8'b00000000 ;
			15'h00005220 : data <= 8'b00000000 ;
			15'h00005221 : data <= 8'b00000000 ;
			15'h00005222 : data <= 8'b00000000 ;
			15'h00005223 : data <= 8'b00000000 ;
			15'h00005224 : data <= 8'b00000000 ;
			15'h00005225 : data <= 8'b00000000 ;
			15'h00005226 : data <= 8'b00000000 ;
			15'h00005227 : data <= 8'b00000000 ;
			15'h00005228 : data <= 8'b00000000 ;
			15'h00005229 : data <= 8'b00000000 ;
			15'h0000522A : data <= 8'b00000000 ;
			15'h0000522B : data <= 8'b00000000 ;
			15'h0000522C : data <= 8'b00000000 ;
			15'h0000522D : data <= 8'b00000000 ;
			15'h0000522E : data <= 8'b00000000 ;
			15'h0000522F : data <= 8'b00000000 ;
			15'h00005230 : data <= 8'b00000000 ;
			15'h00005231 : data <= 8'b00000000 ;
			15'h00005232 : data <= 8'b00000000 ;
			15'h00005233 : data <= 8'b00000000 ;
			15'h00005234 : data <= 8'b00000000 ;
			15'h00005235 : data <= 8'b00000000 ;
			15'h00005236 : data <= 8'b00000000 ;
			15'h00005237 : data <= 8'b00000000 ;
			15'h00005238 : data <= 8'b00000000 ;
			15'h00005239 : data <= 8'b00000000 ;
			15'h0000523A : data <= 8'b00000000 ;
			15'h0000523B : data <= 8'b00000000 ;
			15'h0000523C : data <= 8'b00000000 ;
			15'h0000523D : data <= 8'b00000000 ;
			15'h0000523E : data <= 8'b00000000 ;
			15'h0000523F : data <= 8'b00000000 ;
			15'h00005240 : data <= 8'b00000000 ;
			15'h00005241 : data <= 8'b00000000 ;
			15'h00005242 : data <= 8'b00000000 ;
			15'h00005243 : data <= 8'b00000000 ;
			15'h00005244 : data <= 8'b00000000 ;
			15'h00005245 : data <= 8'b00000000 ;
			15'h00005246 : data <= 8'b00000000 ;
			15'h00005247 : data <= 8'b00000000 ;
			15'h00005248 : data <= 8'b00000000 ;
			15'h00005249 : data <= 8'b00000000 ;
			15'h0000524A : data <= 8'b00000000 ;
			15'h0000524B : data <= 8'b00000000 ;
			15'h0000524C : data <= 8'b00000000 ;
			15'h0000524D : data <= 8'b00000000 ;
			15'h0000524E : data <= 8'b00000000 ;
			15'h0000524F : data <= 8'b00000000 ;
			15'h00005250 : data <= 8'b00000000 ;
			15'h00005251 : data <= 8'b00000000 ;
			15'h00005252 : data <= 8'b00000000 ;
			15'h00005253 : data <= 8'b00000000 ;
			15'h00005254 : data <= 8'b00000000 ;
			15'h00005255 : data <= 8'b00000000 ;
			15'h00005256 : data <= 8'b00000000 ;
			15'h00005257 : data <= 8'b00000000 ;
			15'h00005258 : data <= 8'b00000000 ;
			15'h00005259 : data <= 8'b00000000 ;
			15'h0000525A : data <= 8'b00000000 ;
			15'h0000525B : data <= 8'b00000000 ;
			15'h0000525C : data <= 8'b00000000 ;
			15'h0000525D : data <= 8'b00000000 ;
			15'h0000525E : data <= 8'b00000000 ;
			15'h0000525F : data <= 8'b00000000 ;
			15'h00005260 : data <= 8'b00000000 ;
			15'h00005261 : data <= 8'b00000000 ;
			15'h00005262 : data <= 8'b00000000 ;
			15'h00005263 : data <= 8'b00000000 ;
			15'h00005264 : data <= 8'b00000000 ;
			15'h00005265 : data <= 8'b00000000 ;
			15'h00005266 : data <= 8'b00000000 ;
			15'h00005267 : data <= 8'b00000000 ;
			15'h00005268 : data <= 8'b00000000 ;
			15'h00005269 : data <= 8'b00000000 ;
			15'h0000526A : data <= 8'b00000000 ;
			15'h0000526B : data <= 8'b00000000 ;
			15'h0000526C : data <= 8'b00000000 ;
			15'h0000526D : data <= 8'b00000000 ;
			15'h0000526E : data <= 8'b00000000 ;
			15'h0000526F : data <= 8'b00000000 ;
			15'h00005270 : data <= 8'b00000000 ;
			15'h00005271 : data <= 8'b00000000 ;
			15'h00005272 : data <= 8'b00000000 ;
			15'h00005273 : data <= 8'b00000000 ;
			15'h00005274 : data <= 8'b00000000 ;
			15'h00005275 : data <= 8'b00000000 ;
			15'h00005276 : data <= 8'b00000000 ;
			15'h00005277 : data <= 8'b00000000 ;
			15'h00005278 : data <= 8'b00000000 ;
			15'h00005279 : data <= 8'b00000000 ;
			15'h0000527A : data <= 8'b00000000 ;
			15'h0000527B : data <= 8'b00000000 ;
			15'h0000527C : data <= 8'b00000000 ;
			15'h0000527D : data <= 8'b00000000 ;
			15'h0000527E : data <= 8'b00000000 ;
			15'h0000527F : data <= 8'b00000000 ;
			15'h00005280 : data <= 8'b00000000 ;
			15'h00005281 : data <= 8'b00000000 ;
			15'h00005282 : data <= 8'b00000000 ;
			15'h00005283 : data <= 8'b00000000 ;
			15'h00005284 : data <= 8'b00000000 ;
			15'h00005285 : data <= 8'b00000000 ;
			15'h00005286 : data <= 8'b00000000 ;
			15'h00005287 : data <= 8'b00000000 ;
			15'h00005288 : data <= 8'b00000000 ;
			15'h00005289 : data <= 8'b00000000 ;
			15'h0000528A : data <= 8'b00000000 ;
			15'h0000528B : data <= 8'b00000000 ;
			15'h0000528C : data <= 8'b00000000 ;
			15'h0000528D : data <= 8'b00000000 ;
			15'h0000528E : data <= 8'b00000000 ;
			15'h0000528F : data <= 8'b00000000 ;
			15'h00005290 : data <= 8'b00000000 ;
			15'h00005291 : data <= 8'b00000000 ;
			15'h00005292 : data <= 8'b00000000 ;
			15'h00005293 : data <= 8'b00000000 ;
			15'h00005294 : data <= 8'b00000000 ;
			15'h00005295 : data <= 8'b00000000 ;
			15'h00005296 : data <= 8'b00000000 ;
			15'h00005297 : data <= 8'b00000000 ;
			15'h00005298 : data <= 8'b00000000 ;
			15'h00005299 : data <= 8'b00000000 ;
			15'h0000529A : data <= 8'b00000000 ;
			15'h0000529B : data <= 8'b00000000 ;
			15'h0000529C : data <= 8'b00000000 ;
			15'h0000529D : data <= 8'b00000000 ;
			15'h0000529E : data <= 8'b00000000 ;
			15'h0000529F : data <= 8'b00000000 ;
			15'h000052A0 : data <= 8'b00000000 ;
			15'h000052A1 : data <= 8'b00000000 ;
			15'h000052A2 : data <= 8'b00000000 ;
			15'h000052A3 : data <= 8'b00000000 ;
			15'h000052A4 : data <= 8'b00000000 ;
			15'h000052A5 : data <= 8'b00000000 ;
			15'h000052A6 : data <= 8'b00000000 ;
			15'h000052A7 : data <= 8'b00000000 ;
			15'h000052A8 : data <= 8'b00000000 ;
			15'h000052A9 : data <= 8'b00000000 ;
			15'h000052AA : data <= 8'b00000000 ;
			15'h000052AB : data <= 8'b00000000 ;
			15'h000052AC : data <= 8'b00000000 ;
			15'h000052AD : data <= 8'b00000000 ;
			15'h000052AE : data <= 8'b00000000 ;
			15'h000052AF : data <= 8'b00000000 ;
			15'h000052B0 : data <= 8'b00000000 ;
			15'h000052B1 : data <= 8'b00000000 ;
			15'h000052B2 : data <= 8'b00000000 ;
			15'h000052B3 : data <= 8'b00000000 ;
			15'h000052B4 : data <= 8'b00000000 ;
			15'h000052B5 : data <= 8'b00000000 ;
			15'h000052B6 : data <= 8'b00000000 ;
			15'h000052B7 : data <= 8'b00000000 ;
			15'h000052B8 : data <= 8'b00000000 ;
			15'h000052B9 : data <= 8'b00000000 ;
			15'h000052BA : data <= 8'b00000000 ;
			15'h000052BB : data <= 8'b00000000 ;
			15'h000052BC : data <= 8'b00000000 ;
			15'h000052BD : data <= 8'b00000000 ;
			15'h000052BE : data <= 8'b00000000 ;
			15'h000052BF : data <= 8'b00000000 ;
			15'h000052C0 : data <= 8'b00000000 ;
			15'h000052C1 : data <= 8'b00000000 ;
			15'h000052C2 : data <= 8'b00000000 ;
			15'h000052C3 : data <= 8'b00000000 ;
			15'h000052C4 : data <= 8'b00000000 ;
			15'h000052C5 : data <= 8'b00000000 ;
			15'h000052C6 : data <= 8'b00000000 ;
			15'h000052C7 : data <= 8'b00000000 ;
			15'h000052C8 : data <= 8'b00000000 ;
			15'h000052C9 : data <= 8'b00000000 ;
			15'h000052CA : data <= 8'b00000000 ;
			15'h000052CB : data <= 8'b00000000 ;
			15'h000052CC : data <= 8'b00000000 ;
			15'h000052CD : data <= 8'b00000000 ;
			15'h000052CE : data <= 8'b00000000 ;
			15'h000052CF : data <= 8'b00000000 ;
			15'h000052D0 : data <= 8'b00000000 ;
			15'h000052D1 : data <= 8'b00000000 ;
			15'h000052D2 : data <= 8'b00000000 ;
			15'h000052D3 : data <= 8'b00000000 ;
			15'h000052D4 : data <= 8'b00000000 ;
			15'h000052D5 : data <= 8'b00000000 ;
			15'h000052D6 : data <= 8'b00000000 ;
			15'h000052D7 : data <= 8'b00000000 ;
			15'h000052D8 : data <= 8'b00000000 ;
			15'h000052D9 : data <= 8'b00000000 ;
			15'h000052DA : data <= 8'b00000000 ;
			15'h000052DB : data <= 8'b00000000 ;
			15'h000052DC : data <= 8'b00000000 ;
			15'h000052DD : data <= 8'b00000000 ;
			15'h000052DE : data <= 8'b00000000 ;
			15'h000052DF : data <= 8'b00000000 ;
			15'h000052E0 : data <= 8'b00000000 ;
			15'h000052E1 : data <= 8'b00000000 ;
			15'h000052E2 : data <= 8'b00000000 ;
			15'h000052E3 : data <= 8'b00000000 ;
			15'h000052E4 : data <= 8'b00000000 ;
			15'h000052E5 : data <= 8'b00000000 ;
			15'h000052E6 : data <= 8'b00000000 ;
			15'h000052E7 : data <= 8'b00000000 ;
			15'h000052E8 : data <= 8'b00000000 ;
			15'h000052E9 : data <= 8'b00000000 ;
			15'h000052EA : data <= 8'b00000000 ;
			15'h000052EB : data <= 8'b00000000 ;
			15'h000052EC : data <= 8'b00000000 ;
			15'h000052ED : data <= 8'b00000000 ;
			15'h000052EE : data <= 8'b00000000 ;
			15'h000052EF : data <= 8'b00000000 ;
			15'h000052F0 : data <= 8'b00000000 ;
			15'h000052F1 : data <= 8'b00000000 ;
			15'h000052F2 : data <= 8'b00000000 ;
			15'h000052F3 : data <= 8'b00000000 ;
			15'h000052F4 : data <= 8'b00000000 ;
			15'h000052F5 : data <= 8'b00000000 ;
			15'h000052F6 : data <= 8'b00000000 ;
			15'h000052F7 : data <= 8'b00000000 ;
			15'h000052F8 : data <= 8'b00000000 ;
			15'h000052F9 : data <= 8'b00000000 ;
			15'h000052FA : data <= 8'b00000000 ;
			15'h000052FB : data <= 8'b00000000 ;
			15'h000052FC : data <= 8'b00000000 ;
			15'h000052FD : data <= 8'b00000000 ;
			15'h000052FE : data <= 8'b00000000 ;
			15'h000052FF : data <= 8'b00000000 ;
			15'h00005300 : data <= 8'b00000000 ;
			15'h00005301 : data <= 8'b00000000 ;
			15'h00005302 : data <= 8'b00000000 ;
			15'h00005303 : data <= 8'b00000000 ;
			15'h00005304 : data <= 8'b00000000 ;
			15'h00005305 : data <= 8'b00000000 ;
			15'h00005306 : data <= 8'b00000000 ;
			15'h00005307 : data <= 8'b00000000 ;
			15'h00005308 : data <= 8'b00000000 ;
			15'h00005309 : data <= 8'b00000000 ;
			15'h0000530A : data <= 8'b00000000 ;
			15'h0000530B : data <= 8'b00000000 ;
			15'h0000530C : data <= 8'b00000000 ;
			15'h0000530D : data <= 8'b00000000 ;
			15'h0000530E : data <= 8'b00000000 ;
			15'h0000530F : data <= 8'b00000000 ;
			15'h00005310 : data <= 8'b00000000 ;
			15'h00005311 : data <= 8'b00000000 ;
			15'h00005312 : data <= 8'b00000000 ;
			15'h00005313 : data <= 8'b00000000 ;
			15'h00005314 : data <= 8'b00000000 ;
			15'h00005315 : data <= 8'b00000000 ;
			15'h00005316 : data <= 8'b00000000 ;
			15'h00005317 : data <= 8'b00000000 ;
			15'h00005318 : data <= 8'b00000000 ;
			15'h00005319 : data <= 8'b00000000 ;
			15'h0000531A : data <= 8'b00000000 ;
			15'h0000531B : data <= 8'b00000000 ;
			15'h0000531C : data <= 8'b00000000 ;
			15'h0000531D : data <= 8'b00000000 ;
			15'h0000531E : data <= 8'b00000000 ;
			15'h0000531F : data <= 8'b00000000 ;
			15'h00005320 : data <= 8'b00000000 ;
			15'h00005321 : data <= 8'b00000000 ;
			15'h00005322 : data <= 8'b00000000 ;
			15'h00005323 : data <= 8'b00000000 ;
			15'h00005324 : data <= 8'b00000000 ;
			15'h00005325 : data <= 8'b00000000 ;
			15'h00005326 : data <= 8'b00000000 ;
			15'h00005327 : data <= 8'b00000000 ;
			15'h00005328 : data <= 8'b00000000 ;
			15'h00005329 : data <= 8'b00000000 ;
			15'h0000532A : data <= 8'b00000000 ;
			15'h0000532B : data <= 8'b00000000 ;
			15'h0000532C : data <= 8'b00000000 ;
			15'h0000532D : data <= 8'b00000000 ;
			15'h0000532E : data <= 8'b00000000 ;
			15'h0000532F : data <= 8'b00000000 ;
			15'h00005330 : data <= 8'b00000000 ;
			15'h00005331 : data <= 8'b00000000 ;
			15'h00005332 : data <= 8'b00000000 ;
			15'h00005333 : data <= 8'b00000000 ;
			15'h00005334 : data <= 8'b00000000 ;
			15'h00005335 : data <= 8'b00000000 ;
			15'h00005336 : data <= 8'b00000000 ;
			15'h00005337 : data <= 8'b00000000 ;
			15'h00005338 : data <= 8'b00000000 ;
			15'h00005339 : data <= 8'b00000000 ;
			15'h0000533A : data <= 8'b00000000 ;
			15'h0000533B : data <= 8'b00000000 ;
			15'h0000533C : data <= 8'b00000000 ;
			15'h0000533D : data <= 8'b00000000 ;
			15'h0000533E : data <= 8'b00000000 ;
			15'h0000533F : data <= 8'b00000000 ;
			15'h00005340 : data <= 8'b00000000 ;
			15'h00005341 : data <= 8'b00000000 ;
			15'h00005342 : data <= 8'b00000000 ;
			15'h00005343 : data <= 8'b00000000 ;
			15'h00005344 : data <= 8'b00000000 ;
			15'h00005345 : data <= 8'b00000000 ;
			15'h00005346 : data <= 8'b00000000 ;
			15'h00005347 : data <= 8'b00000000 ;
			15'h00005348 : data <= 8'b00000000 ;
			15'h00005349 : data <= 8'b00000000 ;
			15'h0000534A : data <= 8'b00000000 ;
			15'h0000534B : data <= 8'b00000000 ;
			15'h0000534C : data <= 8'b00000000 ;
			15'h0000534D : data <= 8'b00000000 ;
			15'h0000534E : data <= 8'b00000000 ;
			15'h0000534F : data <= 8'b00000000 ;
			15'h00005350 : data <= 8'b00000000 ;
			15'h00005351 : data <= 8'b00000000 ;
			15'h00005352 : data <= 8'b00000000 ;
			15'h00005353 : data <= 8'b00000000 ;
			15'h00005354 : data <= 8'b00000000 ;
			15'h00005355 : data <= 8'b00000000 ;
			15'h00005356 : data <= 8'b00000000 ;
			15'h00005357 : data <= 8'b00000000 ;
			15'h00005358 : data <= 8'b00000000 ;
			15'h00005359 : data <= 8'b00000000 ;
			15'h0000535A : data <= 8'b00000000 ;
			15'h0000535B : data <= 8'b00000000 ;
			15'h0000535C : data <= 8'b00000000 ;
			15'h0000535D : data <= 8'b00000000 ;
			15'h0000535E : data <= 8'b00000000 ;
			15'h0000535F : data <= 8'b00000000 ;
			15'h00005360 : data <= 8'b00000000 ;
			15'h00005361 : data <= 8'b00000000 ;
			15'h00005362 : data <= 8'b00000000 ;
			15'h00005363 : data <= 8'b00000000 ;
			15'h00005364 : data <= 8'b00000000 ;
			15'h00005365 : data <= 8'b00000000 ;
			15'h00005366 : data <= 8'b00000000 ;
			15'h00005367 : data <= 8'b00000000 ;
			15'h00005368 : data <= 8'b00000000 ;
			15'h00005369 : data <= 8'b00000000 ;
			15'h0000536A : data <= 8'b00000000 ;
			15'h0000536B : data <= 8'b00000000 ;
			15'h0000536C : data <= 8'b00000000 ;
			15'h0000536D : data <= 8'b00000000 ;
			15'h0000536E : data <= 8'b00000000 ;
			15'h0000536F : data <= 8'b00000000 ;
			15'h00005370 : data <= 8'b00000000 ;
			15'h00005371 : data <= 8'b00000000 ;
			15'h00005372 : data <= 8'b00000000 ;
			15'h00005373 : data <= 8'b00000000 ;
			15'h00005374 : data <= 8'b00000000 ;
			15'h00005375 : data <= 8'b00000000 ;
			15'h00005376 : data <= 8'b00000000 ;
			15'h00005377 : data <= 8'b00000000 ;
			15'h00005378 : data <= 8'b00000000 ;
			15'h00005379 : data <= 8'b00000000 ;
			15'h0000537A : data <= 8'b00000000 ;
			15'h0000537B : data <= 8'b00000000 ;
			15'h0000537C : data <= 8'b00000000 ;
			15'h0000537D : data <= 8'b00000000 ;
			15'h0000537E : data <= 8'b00000000 ;
			15'h0000537F : data <= 8'b00000000 ;
			15'h00005380 : data <= 8'b00000000 ;
			15'h00005381 : data <= 8'b00000000 ;
			15'h00005382 : data <= 8'b00000000 ;
			15'h00005383 : data <= 8'b00000000 ;
			15'h00005384 : data <= 8'b00000000 ;
			15'h00005385 : data <= 8'b00000000 ;
			15'h00005386 : data <= 8'b00000000 ;
			15'h00005387 : data <= 8'b00000000 ;
			15'h00005388 : data <= 8'b00000000 ;
			15'h00005389 : data <= 8'b00000000 ;
			15'h0000538A : data <= 8'b00000000 ;
			15'h0000538B : data <= 8'b00000000 ;
			15'h0000538C : data <= 8'b00000000 ;
			15'h0000538D : data <= 8'b00000000 ;
			15'h0000538E : data <= 8'b00000000 ;
			15'h0000538F : data <= 8'b00000000 ;
			15'h00005390 : data <= 8'b00000000 ;
			15'h00005391 : data <= 8'b00000000 ;
			15'h00005392 : data <= 8'b00000000 ;
			15'h00005393 : data <= 8'b00000000 ;
			15'h00005394 : data <= 8'b00000000 ;
			15'h00005395 : data <= 8'b00000000 ;
			15'h00005396 : data <= 8'b00000000 ;
			15'h00005397 : data <= 8'b00000000 ;
			15'h00005398 : data <= 8'b00000000 ;
			15'h00005399 : data <= 8'b00000000 ;
			15'h0000539A : data <= 8'b00000000 ;
			15'h0000539B : data <= 8'b00000000 ;
			15'h0000539C : data <= 8'b00000000 ;
			15'h0000539D : data <= 8'b00000000 ;
			15'h0000539E : data <= 8'b00000000 ;
			15'h0000539F : data <= 8'b00000000 ;
			15'h000053A0 : data <= 8'b00000000 ;
			15'h000053A1 : data <= 8'b00000000 ;
			15'h000053A2 : data <= 8'b00000000 ;
			15'h000053A3 : data <= 8'b00000000 ;
			15'h000053A4 : data <= 8'b00000000 ;
			15'h000053A5 : data <= 8'b00000000 ;
			15'h000053A6 : data <= 8'b00000000 ;
			15'h000053A7 : data <= 8'b00000000 ;
			15'h000053A8 : data <= 8'b00000000 ;
			15'h000053A9 : data <= 8'b00000000 ;
			15'h000053AA : data <= 8'b00000000 ;
			15'h000053AB : data <= 8'b00000000 ;
			15'h000053AC : data <= 8'b00000000 ;
			15'h000053AD : data <= 8'b00000000 ;
			15'h000053AE : data <= 8'b00000000 ;
			15'h000053AF : data <= 8'b00000000 ;
			15'h000053B0 : data <= 8'b00000000 ;
			15'h000053B1 : data <= 8'b00000000 ;
			15'h000053B2 : data <= 8'b00000000 ;
			15'h000053B3 : data <= 8'b00000000 ;
			15'h000053B4 : data <= 8'b00000000 ;
			15'h000053B5 : data <= 8'b00000000 ;
			15'h000053B6 : data <= 8'b00000000 ;
			15'h000053B7 : data <= 8'b00000000 ;
			15'h000053B8 : data <= 8'b00000000 ;
			15'h000053B9 : data <= 8'b00000000 ;
			15'h000053BA : data <= 8'b00000000 ;
			15'h000053BB : data <= 8'b00000000 ;
			15'h000053BC : data <= 8'b00000000 ;
			15'h000053BD : data <= 8'b00000000 ;
			15'h000053BE : data <= 8'b00000000 ;
			15'h000053BF : data <= 8'b00000000 ;
			15'h000053C0 : data <= 8'b00000000 ;
			15'h000053C1 : data <= 8'b00000000 ;
			15'h000053C2 : data <= 8'b00000000 ;
			15'h000053C3 : data <= 8'b00000000 ;
			15'h000053C4 : data <= 8'b00000000 ;
			15'h000053C5 : data <= 8'b00000000 ;
			15'h000053C6 : data <= 8'b00000000 ;
			15'h000053C7 : data <= 8'b00000000 ;
			15'h000053C8 : data <= 8'b00000000 ;
			15'h000053C9 : data <= 8'b00000000 ;
			15'h000053CA : data <= 8'b00000000 ;
			15'h000053CB : data <= 8'b00000000 ;
			15'h000053CC : data <= 8'b00000000 ;
			15'h000053CD : data <= 8'b00000000 ;
			15'h000053CE : data <= 8'b00000000 ;
			15'h000053CF : data <= 8'b00000000 ;
			15'h000053D0 : data <= 8'b00000000 ;
			15'h000053D1 : data <= 8'b00000000 ;
			15'h000053D2 : data <= 8'b00000000 ;
			15'h000053D3 : data <= 8'b00000000 ;
			15'h000053D4 : data <= 8'b00000000 ;
			15'h000053D5 : data <= 8'b00000000 ;
			15'h000053D6 : data <= 8'b00000000 ;
			15'h000053D7 : data <= 8'b00000000 ;
			15'h000053D8 : data <= 8'b00000000 ;
			15'h000053D9 : data <= 8'b00000000 ;
			15'h000053DA : data <= 8'b00000000 ;
			15'h000053DB : data <= 8'b00000000 ;
			15'h000053DC : data <= 8'b00000000 ;
			15'h000053DD : data <= 8'b00000000 ;
			15'h000053DE : data <= 8'b00000000 ;
			15'h000053DF : data <= 8'b00000000 ;
			15'h000053E0 : data <= 8'b00000000 ;
			15'h000053E1 : data <= 8'b00000000 ;
			15'h000053E2 : data <= 8'b00000000 ;
			15'h000053E3 : data <= 8'b00000000 ;
			15'h000053E4 : data <= 8'b00000000 ;
			15'h000053E5 : data <= 8'b00000000 ;
			15'h000053E6 : data <= 8'b00000000 ;
			15'h000053E7 : data <= 8'b00000000 ;
			15'h000053E8 : data <= 8'b00000000 ;
			15'h000053E9 : data <= 8'b00000000 ;
			15'h000053EA : data <= 8'b00000000 ;
			15'h000053EB : data <= 8'b00000000 ;
			15'h000053EC : data <= 8'b00000000 ;
			15'h000053ED : data <= 8'b00000000 ;
			15'h000053EE : data <= 8'b00000000 ;
			15'h000053EF : data <= 8'b00000000 ;
			15'h000053F0 : data <= 8'b00000000 ;
			15'h000053F1 : data <= 8'b00000000 ;
			15'h000053F2 : data <= 8'b00000000 ;
			15'h000053F3 : data <= 8'b00000000 ;
			15'h000053F4 : data <= 8'b00000000 ;
			15'h000053F5 : data <= 8'b00000000 ;
			15'h000053F6 : data <= 8'b00000000 ;
			15'h000053F7 : data <= 8'b00000000 ;
			15'h000053F8 : data <= 8'b00000000 ;
			15'h000053F9 : data <= 8'b00000000 ;
			15'h000053FA : data <= 8'b00000000 ;
			15'h000053FB : data <= 8'b00000000 ;
			15'h000053FC : data <= 8'b00000000 ;
			15'h000053FD : data <= 8'b00000000 ;
			15'h000053FE : data <= 8'b00000000 ;
			15'h000053FF : data <= 8'b00000000 ;
			15'h00005400 : data <= 8'b00000000 ;
			15'h00005401 : data <= 8'b00000000 ;
			15'h00005402 : data <= 8'b00000000 ;
			15'h00005403 : data <= 8'b00000000 ;
			15'h00005404 : data <= 8'b00000000 ;
			15'h00005405 : data <= 8'b00000000 ;
			15'h00005406 : data <= 8'b00000000 ;
			15'h00005407 : data <= 8'b00000000 ;
			15'h00005408 : data <= 8'b00000000 ;
			15'h00005409 : data <= 8'b00000000 ;
			15'h0000540A : data <= 8'b00000000 ;
			15'h0000540B : data <= 8'b00000000 ;
			15'h0000540C : data <= 8'b00000000 ;
			15'h0000540D : data <= 8'b00000000 ;
			15'h0000540E : data <= 8'b00000000 ;
			15'h0000540F : data <= 8'b00000000 ;
			15'h00005410 : data <= 8'b00000000 ;
			15'h00005411 : data <= 8'b00000000 ;
			15'h00005412 : data <= 8'b00000000 ;
			15'h00005413 : data <= 8'b00000000 ;
			15'h00005414 : data <= 8'b00000000 ;
			15'h00005415 : data <= 8'b00000000 ;
			15'h00005416 : data <= 8'b00000000 ;
			15'h00005417 : data <= 8'b00000000 ;
			15'h00005418 : data <= 8'b00000000 ;
			15'h00005419 : data <= 8'b00000000 ;
			15'h0000541A : data <= 8'b00000000 ;
			15'h0000541B : data <= 8'b00000000 ;
			15'h0000541C : data <= 8'b00000000 ;
			15'h0000541D : data <= 8'b00000000 ;
			15'h0000541E : data <= 8'b00000000 ;
			15'h0000541F : data <= 8'b00000000 ;
			15'h00005420 : data <= 8'b00000000 ;
			15'h00005421 : data <= 8'b00000000 ;
			15'h00005422 : data <= 8'b00000000 ;
			15'h00005423 : data <= 8'b00000000 ;
			15'h00005424 : data <= 8'b00000000 ;
			15'h00005425 : data <= 8'b00000000 ;
			15'h00005426 : data <= 8'b00000000 ;
			15'h00005427 : data <= 8'b00000000 ;
			15'h00005428 : data <= 8'b00000000 ;
			15'h00005429 : data <= 8'b00000000 ;
			15'h0000542A : data <= 8'b00000000 ;
			15'h0000542B : data <= 8'b00000000 ;
			15'h0000542C : data <= 8'b00000000 ;
			15'h0000542D : data <= 8'b00000000 ;
			15'h0000542E : data <= 8'b00000000 ;
			15'h0000542F : data <= 8'b00000000 ;
			15'h00005430 : data <= 8'b00000000 ;
			15'h00005431 : data <= 8'b00000000 ;
			15'h00005432 : data <= 8'b00000000 ;
			15'h00005433 : data <= 8'b00000000 ;
			15'h00005434 : data <= 8'b00000000 ;
			15'h00005435 : data <= 8'b00000000 ;
			15'h00005436 : data <= 8'b00000000 ;
			15'h00005437 : data <= 8'b00000000 ;
			15'h00005438 : data <= 8'b00000000 ;
			15'h00005439 : data <= 8'b00000000 ;
			15'h0000543A : data <= 8'b00000000 ;
			15'h0000543B : data <= 8'b00000000 ;
			15'h0000543C : data <= 8'b00000000 ;
			15'h0000543D : data <= 8'b00000000 ;
			15'h0000543E : data <= 8'b00000000 ;
			15'h0000543F : data <= 8'b00000000 ;
			15'h00005440 : data <= 8'b00000000 ;
			15'h00005441 : data <= 8'b00000000 ;
			15'h00005442 : data <= 8'b00000000 ;
			15'h00005443 : data <= 8'b00000000 ;
			15'h00005444 : data <= 8'b00000000 ;
			15'h00005445 : data <= 8'b00000000 ;
			15'h00005446 : data <= 8'b00000000 ;
			15'h00005447 : data <= 8'b00000000 ;
			15'h00005448 : data <= 8'b00000000 ;
			15'h00005449 : data <= 8'b00000000 ;
			15'h0000544A : data <= 8'b00000000 ;
			15'h0000544B : data <= 8'b00000000 ;
			15'h0000544C : data <= 8'b00000000 ;
			15'h0000544D : data <= 8'b00000000 ;
			15'h0000544E : data <= 8'b00000000 ;
			15'h0000544F : data <= 8'b00000000 ;
			15'h00005450 : data <= 8'b00000000 ;
			15'h00005451 : data <= 8'b00000000 ;
			15'h00005452 : data <= 8'b00000000 ;
			15'h00005453 : data <= 8'b00000000 ;
			15'h00005454 : data <= 8'b00000000 ;
			15'h00005455 : data <= 8'b00000000 ;
			15'h00005456 : data <= 8'b00000000 ;
			15'h00005457 : data <= 8'b00000000 ;
			15'h00005458 : data <= 8'b00000000 ;
			15'h00005459 : data <= 8'b00000000 ;
			15'h0000545A : data <= 8'b00000000 ;
			15'h0000545B : data <= 8'b00000000 ;
			15'h0000545C : data <= 8'b00000000 ;
			15'h0000545D : data <= 8'b00000000 ;
			15'h0000545E : data <= 8'b00000000 ;
			15'h0000545F : data <= 8'b00000000 ;
			15'h00005460 : data <= 8'b00000000 ;
			15'h00005461 : data <= 8'b00000000 ;
			15'h00005462 : data <= 8'b00000000 ;
			15'h00005463 : data <= 8'b00000000 ;
			15'h00005464 : data <= 8'b00000000 ;
			15'h00005465 : data <= 8'b00000000 ;
			15'h00005466 : data <= 8'b00000000 ;
			15'h00005467 : data <= 8'b00000000 ;
			15'h00005468 : data <= 8'b00000000 ;
			15'h00005469 : data <= 8'b00000000 ;
			15'h0000546A : data <= 8'b00000000 ;
			15'h0000546B : data <= 8'b00000000 ;
			15'h0000546C : data <= 8'b00000000 ;
			15'h0000546D : data <= 8'b00000000 ;
			15'h0000546E : data <= 8'b00000000 ;
			15'h0000546F : data <= 8'b00000000 ;
			15'h00005470 : data <= 8'b00000000 ;
			15'h00005471 : data <= 8'b00000000 ;
			15'h00005472 : data <= 8'b00000000 ;
			15'h00005473 : data <= 8'b00000000 ;
			15'h00005474 : data <= 8'b00000000 ;
			15'h00005475 : data <= 8'b00000000 ;
			15'h00005476 : data <= 8'b00000000 ;
			15'h00005477 : data <= 8'b00000000 ;
			15'h00005478 : data <= 8'b00000000 ;
			15'h00005479 : data <= 8'b00000000 ;
			15'h0000547A : data <= 8'b00000000 ;
			15'h0000547B : data <= 8'b00000000 ;
			15'h0000547C : data <= 8'b00000000 ;
			15'h0000547D : data <= 8'b00000000 ;
			15'h0000547E : data <= 8'b00000000 ;
			15'h0000547F : data <= 8'b00000000 ;
			15'h00005480 : data <= 8'b00000000 ;
			15'h00005481 : data <= 8'b00000000 ;
			15'h00005482 : data <= 8'b00000000 ;
			15'h00005483 : data <= 8'b00000000 ;
			15'h00005484 : data <= 8'b00000000 ;
			15'h00005485 : data <= 8'b00000000 ;
			15'h00005486 : data <= 8'b00000000 ;
			15'h00005487 : data <= 8'b00000000 ;
			15'h00005488 : data <= 8'b00000000 ;
			15'h00005489 : data <= 8'b00000000 ;
			15'h0000548A : data <= 8'b00000000 ;
			15'h0000548B : data <= 8'b00000000 ;
			15'h0000548C : data <= 8'b00000000 ;
			15'h0000548D : data <= 8'b00000000 ;
			15'h0000548E : data <= 8'b00000000 ;
			15'h0000548F : data <= 8'b00000000 ;
			15'h00005490 : data <= 8'b00000000 ;
			15'h00005491 : data <= 8'b00000000 ;
			15'h00005492 : data <= 8'b00000000 ;
			15'h00005493 : data <= 8'b00000000 ;
			15'h00005494 : data <= 8'b00000000 ;
			15'h00005495 : data <= 8'b00000000 ;
			15'h00005496 : data <= 8'b00000000 ;
			15'h00005497 : data <= 8'b00000000 ;
			15'h00005498 : data <= 8'b00000000 ;
			15'h00005499 : data <= 8'b00000000 ;
			15'h0000549A : data <= 8'b00000000 ;
			15'h0000549B : data <= 8'b00000000 ;
			15'h0000549C : data <= 8'b00000000 ;
			15'h0000549D : data <= 8'b00000000 ;
			15'h0000549E : data <= 8'b00000000 ;
			15'h0000549F : data <= 8'b00000000 ;
			15'h000054A0 : data <= 8'b00000000 ;
			15'h000054A1 : data <= 8'b00000000 ;
			15'h000054A2 : data <= 8'b00000000 ;
			15'h000054A3 : data <= 8'b00000000 ;
			15'h000054A4 : data <= 8'b00000000 ;
			15'h000054A5 : data <= 8'b00000000 ;
			15'h000054A6 : data <= 8'b00000000 ;
			15'h000054A7 : data <= 8'b00000000 ;
			15'h000054A8 : data <= 8'b00000000 ;
			15'h000054A9 : data <= 8'b00000000 ;
			15'h000054AA : data <= 8'b00000000 ;
			15'h000054AB : data <= 8'b00000000 ;
			15'h000054AC : data <= 8'b00000000 ;
			15'h000054AD : data <= 8'b00000000 ;
			15'h000054AE : data <= 8'b00000000 ;
			15'h000054AF : data <= 8'b00000000 ;
			15'h000054B0 : data <= 8'b00000000 ;
			15'h000054B1 : data <= 8'b00000000 ;
			15'h000054B2 : data <= 8'b00000000 ;
			15'h000054B3 : data <= 8'b00000000 ;
			15'h000054B4 : data <= 8'b00000000 ;
			15'h000054B5 : data <= 8'b00000000 ;
			15'h000054B6 : data <= 8'b00000000 ;
			15'h000054B7 : data <= 8'b00000000 ;
			15'h000054B8 : data <= 8'b00000000 ;
			15'h000054B9 : data <= 8'b00000000 ;
			15'h000054BA : data <= 8'b00000000 ;
			15'h000054BB : data <= 8'b00000000 ;
			15'h000054BC : data <= 8'b00000000 ;
			15'h000054BD : data <= 8'b00000000 ;
			15'h000054BE : data <= 8'b00000000 ;
			15'h000054BF : data <= 8'b00000000 ;
			15'h000054C0 : data <= 8'b00000000 ;
			15'h000054C1 : data <= 8'b00000000 ;
			15'h000054C2 : data <= 8'b00000000 ;
			15'h000054C3 : data <= 8'b00000000 ;
			15'h000054C4 : data <= 8'b00000000 ;
			15'h000054C5 : data <= 8'b00000000 ;
			15'h000054C6 : data <= 8'b00000000 ;
			15'h000054C7 : data <= 8'b00000000 ;
			15'h000054C8 : data <= 8'b00000000 ;
			15'h000054C9 : data <= 8'b00000000 ;
			15'h000054CA : data <= 8'b00000000 ;
			15'h000054CB : data <= 8'b00000000 ;
			15'h000054CC : data <= 8'b00000000 ;
			15'h000054CD : data <= 8'b00000000 ;
			15'h000054CE : data <= 8'b00000000 ;
			15'h000054CF : data <= 8'b00000000 ;
			15'h000054D0 : data <= 8'b00000000 ;
			15'h000054D1 : data <= 8'b00000000 ;
			15'h000054D2 : data <= 8'b00000000 ;
			15'h000054D3 : data <= 8'b00000000 ;
			15'h000054D4 : data <= 8'b00000000 ;
			15'h000054D5 : data <= 8'b00000000 ;
			15'h000054D6 : data <= 8'b00000000 ;
			15'h000054D7 : data <= 8'b00000000 ;
			15'h000054D8 : data <= 8'b00000000 ;
			15'h000054D9 : data <= 8'b00000000 ;
			15'h000054DA : data <= 8'b00000000 ;
			15'h000054DB : data <= 8'b00000000 ;
			15'h000054DC : data <= 8'b00000000 ;
			15'h000054DD : data <= 8'b00000000 ;
			15'h000054DE : data <= 8'b00000000 ;
			15'h000054DF : data <= 8'b00000000 ;
			15'h000054E0 : data <= 8'b00000000 ;
			15'h000054E1 : data <= 8'b00000000 ;
			15'h000054E2 : data <= 8'b00000000 ;
			15'h000054E3 : data <= 8'b00000000 ;
			15'h000054E4 : data <= 8'b00000000 ;
			15'h000054E5 : data <= 8'b00000000 ;
			15'h000054E6 : data <= 8'b00000000 ;
			15'h000054E7 : data <= 8'b00000000 ;
			15'h000054E8 : data <= 8'b00000000 ;
			15'h000054E9 : data <= 8'b00000000 ;
			15'h000054EA : data <= 8'b00000000 ;
			15'h000054EB : data <= 8'b00000000 ;
			15'h000054EC : data <= 8'b00000000 ;
			15'h000054ED : data <= 8'b00000000 ;
			15'h000054EE : data <= 8'b00000000 ;
			15'h000054EF : data <= 8'b00000000 ;
			15'h000054F0 : data <= 8'b00000000 ;
			15'h000054F1 : data <= 8'b00000000 ;
			15'h000054F2 : data <= 8'b00000000 ;
			15'h000054F3 : data <= 8'b00000000 ;
			15'h000054F4 : data <= 8'b00000000 ;
			15'h000054F5 : data <= 8'b00000000 ;
			15'h000054F6 : data <= 8'b00000000 ;
			15'h000054F7 : data <= 8'b00000000 ;
			15'h000054F8 : data <= 8'b00000000 ;
			15'h000054F9 : data <= 8'b00000000 ;
			15'h000054FA : data <= 8'b00000000 ;
			15'h000054FB : data <= 8'b00000000 ;
			15'h000054FC : data <= 8'b00000000 ;
			15'h000054FD : data <= 8'b00000000 ;
			15'h000054FE : data <= 8'b00000000 ;
			15'h000054FF : data <= 8'b00000000 ;
			15'h00005500 : data <= 8'b00000000 ;
			15'h00005501 : data <= 8'b00000000 ;
			15'h00005502 : data <= 8'b00000000 ;
			15'h00005503 : data <= 8'b00000000 ;
			15'h00005504 : data <= 8'b00000000 ;
			15'h00005505 : data <= 8'b00000000 ;
			15'h00005506 : data <= 8'b00000000 ;
			15'h00005507 : data <= 8'b00000000 ;
			15'h00005508 : data <= 8'b00000000 ;
			15'h00005509 : data <= 8'b00000000 ;
			15'h0000550A : data <= 8'b00000000 ;
			15'h0000550B : data <= 8'b00000000 ;
			15'h0000550C : data <= 8'b00000000 ;
			15'h0000550D : data <= 8'b00000000 ;
			15'h0000550E : data <= 8'b00000000 ;
			15'h0000550F : data <= 8'b00000000 ;
			15'h00005510 : data <= 8'b00000000 ;
			15'h00005511 : data <= 8'b00000000 ;
			15'h00005512 : data <= 8'b00000000 ;
			15'h00005513 : data <= 8'b00000000 ;
			15'h00005514 : data <= 8'b00000000 ;
			15'h00005515 : data <= 8'b00000000 ;
			15'h00005516 : data <= 8'b00000000 ;
			15'h00005517 : data <= 8'b00000000 ;
			15'h00005518 : data <= 8'b00000000 ;
			15'h00005519 : data <= 8'b00000000 ;
			15'h0000551A : data <= 8'b00000000 ;
			15'h0000551B : data <= 8'b00000000 ;
			15'h0000551C : data <= 8'b00000000 ;
			15'h0000551D : data <= 8'b00000000 ;
			15'h0000551E : data <= 8'b00000000 ;
			15'h0000551F : data <= 8'b00000000 ;
			15'h00005520 : data <= 8'b00000000 ;
			15'h00005521 : data <= 8'b00000000 ;
			15'h00005522 : data <= 8'b00000000 ;
			15'h00005523 : data <= 8'b00000000 ;
			15'h00005524 : data <= 8'b00000000 ;
			15'h00005525 : data <= 8'b00000000 ;
			15'h00005526 : data <= 8'b00000000 ;
			15'h00005527 : data <= 8'b00000000 ;
			15'h00005528 : data <= 8'b00000000 ;
			15'h00005529 : data <= 8'b00000000 ;
			15'h0000552A : data <= 8'b00000000 ;
			15'h0000552B : data <= 8'b00000000 ;
			15'h0000552C : data <= 8'b00000000 ;
			15'h0000552D : data <= 8'b00000000 ;
			15'h0000552E : data <= 8'b00000000 ;
			15'h0000552F : data <= 8'b00000000 ;
			15'h00005530 : data <= 8'b00000000 ;
			15'h00005531 : data <= 8'b00000000 ;
			15'h00005532 : data <= 8'b00000000 ;
			15'h00005533 : data <= 8'b00000000 ;
			15'h00005534 : data <= 8'b00000000 ;
			15'h00005535 : data <= 8'b00000000 ;
			15'h00005536 : data <= 8'b00000000 ;
			15'h00005537 : data <= 8'b00000000 ;
			15'h00005538 : data <= 8'b00000000 ;
			15'h00005539 : data <= 8'b00000000 ;
			15'h0000553A : data <= 8'b00000000 ;
			15'h0000553B : data <= 8'b00000000 ;
			15'h0000553C : data <= 8'b00000000 ;
			15'h0000553D : data <= 8'b00000000 ;
			15'h0000553E : data <= 8'b00000000 ;
			15'h0000553F : data <= 8'b00000000 ;
			15'h00005540 : data <= 8'b00000000 ;
			15'h00005541 : data <= 8'b00000000 ;
			15'h00005542 : data <= 8'b00000000 ;
			15'h00005543 : data <= 8'b00000000 ;
			15'h00005544 : data <= 8'b00000000 ;
			15'h00005545 : data <= 8'b00000000 ;
			15'h00005546 : data <= 8'b00000000 ;
			15'h00005547 : data <= 8'b00000000 ;
			15'h00005548 : data <= 8'b00000000 ;
			15'h00005549 : data <= 8'b00000000 ;
			15'h0000554A : data <= 8'b00000000 ;
			15'h0000554B : data <= 8'b00000000 ;
			15'h0000554C : data <= 8'b00000000 ;
			15'h0000554D : data <= 8'b00000000 ;
			15'h0000554E : data <= 8'b00000000 ;
			15'h0000554F : data <= 8'b00000000 ;
			15'h00005550 : data <= 8'b00000000 ;
			15'h00005551 : data <= 8'b00000000 ;
			15'h00005552 : data <= 8'b00000000 ;
			15'h00005553 : data <= 8'b00000000 ;
			15'h00005554 : data <= 8'b00000000 ;
			15'h00005555 : data <= 8'b00000000 ;
			15'h00005556 : data <= 8'b00000000 ;
			15'h00005557 : data <= 8'b00000000 ;
			15'h00005558 : data <= 8'b00000000 ;
			15'h00005559 : data <= 8'b00000000 ;
			15'h0000555A : data <= 8'b00000000 ;
			15'h0000555B : data <= 8'b00000000 ;
			15'h0000555C : data <= 8'b00000000 ;
			15'h0000555D : data <= 8'b00000000 ;
			15'h0000555E : data <= 8'b00000000 ;
			15'h0000555F : data <= 8'b00000000 ;
			15'h00005560 : data <= 8'b00000000 ;
			15'h00005561 : data <= 8'b00000000 ;
			15'h00005562 : data <= 8'b00000000 ;
			15'h00005563 : data <= 8'b00000000 ;
			15'h00005564 : data <= 8'b00000000 ;
			15'h00005565 : data <= 8'b00000000 ;
			15'h00005566 : data <= 8'b00000000 ;
			15'h00005567 : data <= 8'b00000000 ;
			15'h00005568 : data <= 8'b00000000 ;
			15'h00005569 : data <= 8'b00000000 ;
			15'h0000556A : data <= 8'b00000000 ;
			15'h0000556B : data <= 8'b00000000 ;
			15'h0000556C : data <= 8'b00000000 ;
			15'h0000556D : data <= 8'b00000000 ;
			15'h0000556E : data <= 8'b00000000 ;
			15'h0000556F : data <= 8'b00000000 ;
			15'h00005570 : data <= 8'b00000000 ;
			15'h00005571 : data <= 8'b00000000 ;
			15'h00005572 : data <= 8'b00000000 ;
			15'h00005573 : data <= 8'b00000000 ;
			15'h00005574 : data <= 8'b00000000 ;
			15'h00005575 : data <= 8'b00000000 ;
			15'h00005576 : data <= 8'b00000000 ;
			15'h00005577 : data <= 8'b00000000 ;
			15'h00005578 : data <= 8'b00000000 ;
			15'h00005579 : data <= 8'b00000000 ;
			15'h0000557A : data <= 8'b00000000 ;
			15'h0000557B : data <= 8'b00000000 ;
			15'h0000557C : data <= 8'b00000000 ;
			15'h0000557D : data <= 8'b00000000 ;
			15'h0000557E : data <= 8'b00000000 ;
			15'h0000557F : data <= 8'b00000000 ;
			15'h00005580 : data <= 8'b00000000 ;
			15'h00005581 : data <= 8'b00000000 ;
			15'h00005582 : data <= 8'b00000000 ;
			15'h00005583 : data <= 8'b00000000 ;
			15'h00005584 : data <= 8'b00000000 ;
			15'h00005585 : data <= 8'b00000000 ;
			15'h00005586 : data <= 8'b00000000 ;
			15'h00005587 : data <= 8'b00000000 ;
			15'h00005588 : data <= 8'b00000000 ;
			15'h00005589 : data <= 8'b00000000 ;
			15'h0000558A : data <= 8'b00000000 ;
			15'h0000558B : data <= 8'b00000000 ;
			15'h0000558C : data <= 8'b00000000 ;
			15'h0000558D : data <= 8'b00000000 ;
			15'h0000558E : data <= 8'b00000000 ;
			15'h0000558F : data <= 8'b00000000 ;
			15'h00005590 : data <= 8'b00000000 ;
			15'h00005591 : data <= 8'b00000000 ;
			15'h00005592 : data <= 8'b00000000 ;
			15'h00005593 : data <= 8'b00000000 ;
			15'h00005594 : data <= 8'b00000000 ;
			15'h00005595 : data <= 8'b00000000 ;
			15'h00005596 : data <= 8'b00000000 ;
			15'h00005597 : data <= 8'b00000000 ;
			15'h00005598 : data <= 8'b00000000 ;
			15'h00005599 : data <= 8'b00000000 ;
			15'h0000559A : data <= 8'b00000000 ;
			15'h0000559B : data <= 8'b00000000 ;
			15'h0000559C : data <= 8'b00000000 ;
			15'h0000559D : data <= 8'b00000000 ;
			15'h0000559E : data <= 8'b00000000 ;
			15'h0000559F : data <= 8'b00000000 ;
			15'h000055A0 : data <= 8'b00000000 ;
			15'h000055A1 : data <= 8'b00000000 ;
			15'h000055A2 : data <= 8'b00000000 ;
			15'h000055A3 : data <= 8'b00000000 ;
			15'h000055A4 : data <= 8'b00000000 ;
			15'h000055A5 : data <= 8'b00000000 ;
			15'h000055A6 : data <= 8'b00000000 ;
			15'h000055A7 : data <= 8'b00000000 ;
			15'h000055A8 : data <= 8'b00000000 ;
			15'h000055A9 : data <= 8'b00000000 ;
			15'h000055AA : data <= 8'b00000000 ;
			15'h000055AB : data <= 8'b00000000 ;
			15'h000055AC : data <= 8'b00000000 ;
			15'h000055AD : data <= 8'b00000000 ;
			15'h000055AE : data <= 8'b00000000 ;
			15'h000055AF : data <= 8'b00000000 ;
			15'h000055B0 : data <= 8'b00000000 ;
			15'h000055B1 : data <= 8'b00000000 ;
			15'h000055B2 : data <= 8'b00000000 ;
			15'h000055B3 : data <= 8'b00000000 ;
			15'h000055B4 : data <= 8'b00000000 ;
			15'h000055B5 : data <= 8'b00000000 ;
			15'h000055B6 : data <= 8'b00000000 ;
			15'h000055B7 : data <= 8'b00000000 ;
			15'h000055B8 : data <= 8'b00000000 ;
			15'h000055B9 : data <= 8'b00000000 ;
			15'h000055BA : data <= 8'b00000000 ;
			15'h000055BB : data <= 8'b00000000 ;
			15'h000055BC : data <= 8'b00000000 ;
			15'h000055BD : data <= 8'b00000000 ;
			15'h000055BE : data <= 8'b00000000 ;
			15'h000055BF : data <= 8'b00000000 ;
			15'h000055C0 : data <= 8'b00000000 ;
			15'h000055C1 : data <= 8'b00000000 ;
			15'h000055C2 : data <= 8'b00000000 ;
			15'h000055C3 : data <= 8'b00000000 ;
			15'h000055C4 : data <= 8'b00000000 ;
			15'h000055C5 : data <= 8'b00000000 ;
			15'h000055C6 : data <= 8'b00000000 ;
			15'h000055C7 : data <= 8'b00000000 ;
			15'h000055C8 : data <= 8'b00000000 ;
			15'h000055C9 : data <= 8'b00000000 ;
			15'h000055CA : data <= 8'b00000000 ;
			15'h000055CB : data <= 8'b00000000 ;
			15'h000055CC : data <= 8'b00000000 ;
			15'h000055CD : data <= 8'b00000000 ;
			15'h000055CE : data <= 8'b00000000 ;
			15'h000055CF : data <= 8'b00000000 ;
			15'h000055D0 : data <= 8'b00000000 ;
			15'h000055D1 : data <= 8'b00000000 ;
			15'h000055D2 : data <= 8'b00000000 ;
			15'h000055D3 : data <= 8'b00000000 ;
			15'h000055D4 : data <= 8'b00000000 ;
			15'h000055D5 : data <= 8'b00000000 ;
			15'h000055D6 : data <= 8'b00000000 ;
			15'h000055D7 : data <= 8'b00000000 ;
			15'h000055D8 : data <= 8'b00000000 ;
			15'h000055D9 : data <= 8'b00000000 ;
			15'h000055DA : data <= 8'b00000000 ;
			15'h000055DB : data <= 8'b00000000 ;
			15'h000055DC : data <= 8'b00000000 ;
			15'h000055DD : data <= 8'b00000000 ;
			15'h000055DE : data <= 8'b00000000 ;
			15'h000055DF : data <= 8'b00000000 ;
			15'h000055E0 : data <= 8'b00000000 ;
			15'h000055E1 : data <= 8'b00000000 ;
			15'h000055E2 : data <= 8'b00000000 ;
			15'h000055E3 : data <= 8'b00000000 ;
			15'h000055E4 : data <= 8'b00000000 ;
			15'h000055E5 : data <= 8'b00000000 ;
			15'h000055E6 : data <= 8'b00000000 ;
			15'h000055E7 : data <= 8'b00000000 ;
			15'h000055E8 : data <= 8'b00000000 ;
			15'h000055E9 : data <= 8'b00000000 ;
			15'h000055EA : data <= 8'b00000000 ;
			15'h000055EB : data <= 8'b00000000 ;
			15'h000055EC : data <= 8'b00000000 ;
			15'h000055ED : data <= 8'b00000000 ;
			15'h000055EE : data <= 8'b00000000 ;
			15'h000055EF : data <= 8'b00000000 ;
			15'h000055F0 : data <= 8'b00000000 ;
			15'h000055F1 : data <= 8'b00000000 ;
			15'h000055F2 : data <= 8'b00000000 ;
			15'h000055F3 : data <= 8'b00000000 ;
			15'h000055F4 : data <= 8'b00000000 ;
			15'h000055F5 : data <= 8'b00000000 ;
			15'h000055F6 : data <= 8'b00000000 ;
			15'h000055F7 : data <= 8'b00000000 ;
			15'h000055F8 : data <= 8'b00000000 ;
			15'h000055F9 : data <= 8'b00000000 ;
			15'h000055FA : data <= 8'b00000000 ;
			15'h000055FB : data <= 8'b00000000 ;
			15'h000055FC : data <= 8'b00000000 ;
			15'h000055FD : data <= 8'b00000000 ;
			15'h000055FE : data <= 8'b00000000 ;
			15'h000055FF : data <= 8'b00000000 ;
			15'h00005600 : data <= 8'b00000000 ;
			15'h00005601 : data <= 8'b00000000 ;
			15'h00005602 : data <= 8'b00000000 ;
			15'h00005603 : data <= 8'b00000000 ;
			15'h00005604 : data <= 8'b00000000 ;
			15'h00005605 : data <= 8'b00000000 ;
			15'h00005606 : data <= 8'b00000000 ;
			15'h00005607 : data <= 8'b00000000 ;
			15'h00005608 : data <= 8'b00000000 ;
			15'h00005609 : data <= 8'b00000000 ;
			15'h0000560A : data <= 8'b00000000 ;
			15'h0000560B : data <= 8'b00000000 ;
			15'h0000560C : data <= 8'b00000000 ;
			15'h0000560D : data <= 8'b00000000 ;
			15'h0000560E : data <= 8'b00000000 ;
			15'h0000560F : data <= 8'b00000000 ;
			15'h00005610 : data <= 8'b00000000 ;
			15'h00005611 : data <= 8'b00000000 ;
			15'h00005612 : data <= 8'b00000000 ;
			15'h00005613 : data <= 8'b00000000 ;
			15'h00005614 : data <= 8'b00000000 ;
			15'h00005615 : data <= 8'b00000000 ;
			15'h00005616 : data <= 8'b00000000 ;
			15'h00005617 : data <= 8'b00000000 ;
			15'h00005618 : data <= 8'b00000000 ;
			15'h00005619 : data <= 8'b00000000 ;
			15'h0000561A : data <= 8'b00000000 ;
			15'h0000561B : data <= 8'b00000000 ;
			15'h0000561C : data <= 8'b00000000 ;
			15'h0000561D : data <= 8'b00000000 ;
			15'h0000561E : data <= 8'b00000000 ;
			15'h0000561F : data <= 8'b00000000 ;
			15'h00005620 : data <= 8'b00000000 ;
			15'h00005621 : data <= 8'b00000000 ;
			15'h00005622 : data <= 8'b00000000 ;
			15'h00005623 : data <= 8'b00000000 ;
			15'h00005624 : data <= 8'b00000000 ;
			15'h00005625 : data <= 8'b00000000 ;
			15'h00005626 : data <= 8'b00000000 ;
			15'h00005627 : data <= 8'b00000000 ;
			15'h00005628 : data <= 8'b00000000 ;
			15'h00005629 : data <= 8'b00000000 ;
			15'h0000562A : data <= 8'b00000000 ;
			15'h0000562B : data <= 8'b00000000 ;
			15'h0000562C : data <= 8'b00000000 ;
			15'h0000562D : data <= 8'b00000000 ;
			15'h0000562E : data <= 8'b00000000 ;
			15'h0000562F : data <= 8'b00000000 ;
			15'h00005630 : data <= 8'b00000000 ;
			15'h00005631 : data <= 8'b00000000 ;
			15'h00005632 : data <= 8'b00000000 ;
			15'h00005633 : data <= 8'b00000000 ;
			15'h00005634 : data <= 8'b00000000 ;
			15'h00005635 : data <= 8'b00000000 ;
			15'h00005636 : data <= 8'b00000000 ;
			15'h00005637 : data <= 8'b00000000 ;
			15'h00005638 : data <= 8'b00000000 ;
			15'h00005639 : data <= 8'b00000000 ;
			15'h0000563A : data <= 8'b00000000 ;
			15'h0000563B : data <= 8'b00000000 ;
			15'h0000563C : data <= 8'b00000000 ;
			15'h0000563D : data <= 8'b00000000 ;
			15'h0000563E : data <= 8'b00000000 ;
			15'h0000563F : data <= 8'b00000000 ;
			15'h00005640 : data <= 8'b00000000 ;
			15'h00005641 : data <= 8'b00000000 ;
			15'h00005642 : data <= 8'b00000000 ;
			15'h00005643 : data <= 8'b00000000 ;
			15'h00005644 : data <= 8'b00000000 ;
			15'h00005645 : data <= 8'b00000000 ;
			15'h00005646 : data <= 8'b00000000 ;
			15'h00005647 : data <= 8'b00000000 ;
			15'h00005648 : data <= 8'b00000000 ;
			15'h00005649 : data <= 8'b00000000 ;
			15'h0000564A : data <= 8'b00000000 ;
			15'h0000564B : data <= 8'b00000000 ;
			15'h0000564C : data <= 8'b00000000 ;
			15'h0000564D : data <= 8'b00000000 ;
			15'h0000564E : data <= 8'b00000000 ;
			15'h0000564F : data <= 8'b00000000 ;
			15'h00005650 : data <= 8'b00000000 ;
			15'h00005651 : data <= 8'b00000000 ;
			15'h00005652 : data <= 8'b00000000 ;
			15'h00005653 : data <= 8'b00000000 ;
			15'h00005654 : data <= 8'b00000000 ;
			15'h00005655 : data <= 8'b00000000 ;
			15'h00005656 : data <= 8'b00000000 ;
			15'h00005657 : data <= 8'b00000000 ;
			15'h00005658 : data <= 8'b00000000 ;
			15'h00005659 : data <= 8'b00000000 ;
			15'h0000565A : data <= 8'b00000000 ;
			15'h0000565B : data <= 8'b00000000 ;
			15'h0000565C : data <= 8'b00000000 ;
			15'h0000565D : data <= 8'b00000000 ;
			15'h0000565E : data <= 8'b00000000 ;
			15'h0000565F : data <= 8'b00000000 ;
			15'h00005660 : data <= 8'b00000000 ;
			15'h00005661 : data <= 8'b00000000 ;
			15'h00005662 : data <= 8'b00000000 ;
			15'h00005663 : data <= 8'b00000000 ;
			15'h00005664 : data <= 8'b00000000 ;
			15'h00005665 : data <= 8'b00000000 ;
			15'h00005666 : data <= 8'b00000000 ;
			15'h00005667 : data <= 8'b00000000 ;
			15'h00005668 : data <= 8'b00000000 ;
			15'h00005669 : data <= 8'b00000000 ;
			15'h0000566A : data <= 8'b00000000 ;
			15'h0000566B : data <= 8'b00000000 ;
			15'h0000566C : data <= 8'b00000000 ;
			15'h0000566D : data <= 8'b00000000 ;
			15'h0000566E : data <= 8'b00000000 ;
			15'h0000566F : data <= 8'b00000000 ;
			15'h00005670 : data <= 8'b00000000 ;
			15'h00005671 : data <= 8'b00000000 ;
			15'h00005672 : data <= 8'b00000000 ;
			15'h00005673 : data <= 8'b00000000 ;
			15'h00005674 : data <= 8'b00000000 ;
			15'h00005675 : data <= 8'b00000000 ;
			15'h00005676 : data <= 8'b00000000 ;
			15'h00005677 : data <= 8'b00000000 ;
			15'h00005678 : data <= 8'b00000000 ;
			15'h00005679 : data <= 8'b00000000 ;
			15'h0000567A : data <= 8'b00000000 ;
			15'h0000567B : data <= 8'b00000000 ;
			15'h0000567C : data <= 8'b00000000 ;
			15'h0000567D : data <= 8'b00000000 ;
			15'h0000567E : data <= 8'b00000000 ;
			15'h0000567F : data <= 8'b00000000 ;
			15'h00005680 : data <= 8'b00000000 ;
			15'h00005681 : data <= 8'b00000000 ;
			15'h00005682 : data <= 8'b00000000 ;
			15'h00005683 : data <= 8'b00000000 ;
			15'h00005684 : data <= 8'b00000000 ;
			15'h00005685 : data <= 8'b00000000 ;
			15'h00005686 : data <= 8'b00000000 ;
			15'h00005687 : data <= 8'b00000000 ;
			15'h00005688 : data <= 8'b00000000 ;
			15'h00005689 : data <= 8'b00000000 ;
			15'h0000568A : data <= 8'b00000000 ;
			15'h0000568B : data <= 8'b00000000 ;
			15'h0000568C : data <= 8'b00000000 ;
			15'h0000568D : data <= 8'b00000000 ;
			15'h0000568E : data <= 8'b00000000 ;
			15'h0000568F : data <= 8'b00000000 ;
			15'h00005690 : data <= 8'b00000000 ;
			15'h00005691 : data <= 8'b00000000 ;
			15'h00005692 : data <= 8'b00000000 ;
			15'h00005693 : data <= 8'b00000000 ;
			15'h00005694 : data <= 8'b00000000 ;
			15'h00005695 : data <= 8'b00000000 ;
			15'h00005696 : data <= 8'b00000000 ;
			15'h00005697 : data <= 8'b00000000 ;
			15'h00005698 : data <= 8'b00000000 ;
			15'h00005699 : data <= 8'b00000000 ;
			15'h0000569A : data <= 8'b00000000 ;
			15'h0000569B : data <= 8'b00000000 ;
			15'h0000569C : data <= 8'b00000000 ;
			15'h0000569D : data <= 8'b00000000 ;
			15'h0000569E : data <= 8'b00000000 ;
			15'h0000569F : data <= 8'b00000000 ;
			15'h000056A0 : data <= 8'b00000000 ;
			15'h000056A1 : data <= 8'b00000000 ;
			15'h000056A2 : data <= 8'b00000000 ;
			15'h000056A3 : data <= 8'b00000000 ;
			15'h000056A4 : data <= 8'b00000000 ;
			15'h000056A5 : data <= 8'b00000000 ;
			15'h000056A6 : data <= 8'b00000000 ;
			15'h000056A7 : data <= 8'b00000000 ;
			15'h000056A8 : data <= 8'b00000000 ;
			15'h000056A9 : data <= 8'b00000000 ;
			15'h000056AA : data <= 8'b00000000 ;
			15'h000056AB : data <= 8'b00000000 ;
			15'h000056AC : data <= 8'b00000000 ;
			15'h000056AD : data <= 8'b00000000 ;
			15'h000056AE : data <= 8'b00000000 ;
			15'h000056AF : data <= 8'b00000000 ;
			15'h000056B0 : data <= 8'b00000000 ;
			15'h000056B1 : data <= 8'b00000000 ;
			15'h000056B2 : data <= 8'b00000000 ;
			15'h000056B3 : data <= 8'b00000000 ;
			15'h000056B4 : data <= 8'b00000000 ;
			15'h000056B5 : data <= 8'b00000000 ;
			15'h000056B6 : data <= 8'b00000000 ;
			15'h000056B7 : data <= 8'b00000000 ;
			15'h000056B8 : data <= 8'b00000000 ;
			15'h000056B9 : data <= 8'b00000000 ;
			15'h000056BA : data <= 8'b00000000 ;
			15'h000056BB : data <= 8'b00000000 ;
			15'h000056BC : data <= 8'b00000000 ;
			15'h000056BD : data <= 8'b00000000 ;
			15'h000056BE : data <= 8'b00000000 ;
			15'h000056BF : data <= 8'b00000000 ;
			15'h000056C0 : data <= 8'b00000000 ;
			15'h000056C1 : data <= 8'b00000000 ;
			15'h000056C2 : data <= 8'b00000000 ;
			15'h000056C3 : data <= 8'b00000000 ;
			15'h000056C4 : data <= 8'b00000000 ;
			15'h000056C5 : data <= 8'b00000000 ;
			15'h000056C6 : data <= 8'b00000000 ;
			15'h000056C7 : data <= 8'b00000000 ;
			15'h000056C8 : data <= 8'b00000000 ;
			15'h000056C9 : data <= 8'b00000000 ;
			15'h000056CA : data <= 8'b00000000 ;
			15'h000056CB : data <= 8'b00000000 ;
			15'h000056CC : data <= 8'b00000000 ;
			15'h000056CD : data <= 8'b00000000 ;
			15'h000056CE : data <= 8'b00000000 ;
			15'h000056CF : data <= 8'b00000000 ;
			15'h000056D0 : data <= 8'b00000000 ;
			15'h000056D1 : data <= 8'b00000000 ;
			15'h000056D2 : data <= 8'b00000000 ;
			15'h000056D3 : data <= 8'b00000000 ;
			15'h000056D4 : data <= 8'b00000000 ;
			15'h000056D5 : data <= 8'b00000000 ;
			15'h000056D6 : data <= 8'b00000000 ;
			15'h000056D7 : data <= 8'b00000000 ;
			15'h000056D8 : data <= 8'b00000000 ;
			15'h000056D9 : data <= 8'b00000000 ;
			15'h000056DA : data <= 8'b00000000 ;
			15'h000056DB : data <= 8'b00000000 ;
			15'h000056DC : data <= 8'b00000000 ;
			15'h000056DD : data <= 8'b00000000 ;
			15'h000056DE : data <= 8'b00000000 ;
			15'h000056DF : data <= 8'b00000000 ;
			15'h000056E0 : data <= 8'b00000000 ;
			15'h000056E1 : data <= 8'b00000000 ;
			15'h000056E2 : data <= 8'b00000000 ;
			15'h000056E3 : data <= 8'b00000000 ;
			15'h000056E4 : data <= 8'b00000000 ;
			15'h000056E5 : data <= 8'b00000000 ;
			15'h000056E6 : data <= 8'b00000000 ;
			15'h000056E7 : data <= 8'b00000000 ;
			15'h000056E8 : data <= 8'b00000000 ;
			15'h000056E9 : data <= 8'b00000000 ;
			15'h000056EA : data <= 8'b00000000 ;
			15'h000056EB : data <= 8'b00000000 ;
			15'h000056EC : data <= 8'b00000000 ;
			15'h000056ED : data <= 8'b00000000 ;
			15'h000056EE : data <= 8'b00000000 ;
			15'h000056EF : data <= 8'b00000000 ;
			15'h000056F0 : data <= 8'b00000000 ;
			15'h000056F1 : data <= 8'b00000000 ;
			15'h000056F2 : data <= 8'b00000000 ;
			15'h000056F3 : data <= 8'b00000000 ;
			15'h000056F4 : data <= 8'b00000000 ;
			15'h000056F5 : data <= 8'b00000000 ;
			15'h000056F6 : data <= 8'b00000000 ;
			15'h000056F7 : data <= 8'b00000000 ;
			15'h000056F8 : data <= 8'b00000000 ;
			15'h000056F9 : data <= 8'b00000000 ;
			15'h000056FA : data <= 8'b00000000 ;
			15'h000056FB : data <= 8'b00000000 ;
			15'h000056FC : data <= 8'b00000000 ;
			15'h000056FD : data <= 8'b00000000 ;
			15'h000056FE : data <= 8'b00000000 ;
			15'h000056FF : data <= 8'b00000000 ;
			15'h00005700 : data <= 8'b00000000 ;
			15'h00005701 : data <= 8'b00000000 ;
			15'h00005702 : data <= 8'b00000000 ;
			15'h00005703 : data <= 8'b00000000 ;
			15'h00005704 : data <= 8'b00000000 ;
			15'h00005705 : data <= 8'b00000000 ;
			15'h00005706 : data <= 8'b00000000 ;
			15'h00005707 : data <= 8'b00000000 ;
			15'h00005708 : data <= 8'b00000000 ;
			15'h00005709 : data <= 8'b00000000 ;
			15'h0000570A : data <= 8'b00000000 ;
			15'h0000570B : data <= 8'b00000000 ;
			15'h0000570C : data <= 8'b00000000 ;
			15'h0000570D : data <= 8'b00000000 ;
			15'h0000570E : data <= 8'b00000000 ;
			15'h0000570F : data <= 8'b00000000 ;
			15'h00005710 : data <= 8'b00000000 ;
			15'h00005711 : data <= 8'b00000000 ;
			15'h00005712 : data <= 8'b00000000 ;
			15'h00005713 : data <= 8'b00000000 ;
			15'h00005714 : data <= 8'b00000000 ;
			15'h00005715 : data <= 8'b00000000 ;
			15'h00005716 : data <= 8'b00000000 ;
			15'h00005717 : data <= 8'b00000000 ;
			15'h00005718 : data <= 8'b00000000 ;
			15'h00005719 : data <= 8'b00000000 ;
			15'h0000571A : data <= 8'b00000000 ;
			15'h0000571B : data <= 8'b00000000 ;
			15'h0000571C : data <= 8'b00000000 ;
			15'h0000571D : data <= 8'b00000000 ;
			15'h0000571E : data <= 8'b00000000 ;
			15'h0000571F : data <= 8'b00000000 ;
			15'h00005720 : data <= 8'b00000000 ;
			15'h00005721 : data <= 8'b00000000 ;
			15'h00005722 : data <= 8'b00000000 ;
			15'h00005723 : data <= 8'b00000000 ;
			15'h00005724 : data <= 8'b00000000 ;
			15'h00005725 : data <= 8'b00000000 ;
			15'h00005726 : data <= 8'b00000000 ;
			15'h00005727 : data <= 8'b00000000 ;
			15'h00005728 : data <= 8'b00000000 ;
			15'h00005729 : data <= 8'b00000000 ;
			15'h0000572A : data <= 8'b00000000 ;
			15'h0000572B : data <= 8'b00000000 ;
			15'h0000572C : data <= 8'b00000000 ;
			15'h0000572D : data <= 8'b00000000 ;
			15'h0000572E : data <= 8'b00000000 ;
			15'h0000572F : data <= 8'b00000000 ;
			15'h00005730 : data <= 8'b00000000 ;
			15'h00005731 : data <= 8'b00000000 ;
			15'h00005732 : data <= 8'b00000000 ;
			15'h00005733 : data <= 8'b00000000 ;
			15'h00005734 : data <= 8'b00000000 ;
			15'h00005735 : data <= 8'b00000000 ;
			15'h00005736 : data <= 8'b00000000 ;
			15'h00005737 : data <= 8'b00000000 ;
			15'h00005738 : data <= 8'b00000000 ;
			15'h00005739 : data <= 8'b00000000 ;
			15'h0000573A : data <= 8'b00000000 ;
			15'h0000573B : data <= 8'b00000000 ;
			15'h0000573C : data <= 8'b00000000 ;
			15'h0000573D : data <= 8'b00000000 ;
			15'h0000573E : data <= 8'b00000000 ;
			15'h0000573F : data <= 8'b00000000 ;
			15'h00005740 : data <= 8'b00000000 ;
			15'h00005741 : data <= 8'b00000000 ;
			15'h00005742 : data <= 8'b00000000 ;
			15'h00005743 : data <= 8'b00000000 ;
			15'h00005744 : data <= 8'b00000000 ;
			15'h00005745 : data <= 8'b00000000 ;
			15'h00005746 : data <= 8'b00000000 ;
			15'h00005747 : data <= 8'b00000000 ;
			15'h00005748 : data <= 8'b00000000 ;
			15'h00005749 : data <= 8'b00000000 ;
			15'h0000574A : data <= 8'b00000000 ;
			15'h0000574B : data <= 8'b00000000 ;
			15'h0000574C : data <= 8'b00000000 ;
			15'h0000574D : data <= 8'b00000000 ;
			15'h0000574E : data <= 8'b00000000 ;
			15'h0000574F : data <= 8'b00000000 ;
			15'h00005750 : data <= 8'b00000000 ;
			15'h00005751 : data <= 8'b00000000 ;
			15'h00005752 : data <= 8'b00000000 ;
			15'h00005753 : data <= 8'b00000000 ;
			15'h00005754 : data <= 8'b00000000 ;
			15'h00005755 : data <= 8'b00000000 ;
			15'h00005756 : data <= 8'b00000000 ;
			15'h00005757 : data <= 8'b00000000 ;
			15'h00005758 : data <= 8'b00000000 ;
			15'h00005759 : data <= 8'b00000000 ;
			15'h0000575A : data <= 8'b00000000 ;
			15'h0000575B : data <= 8'b00000000 ;
			15'h0000575C : data <= 8'b00000000 ;
			15'h0000575D : data <= 8'b00000000 ;
			15'h0000575E : data <= 8'b00000000 ;
			15'h0000575F : data <= 8'b00000000 ;
			15'h00005760 : data <= 8'b00000000 ;
			15'h00005761 : data <= 8'b00000000 ;
			15'h00005762 : data <= 8'b00000000 ;
			15'h00005763 : data <= 8'b00000000 ;
			15'h00005764 : data <= 8'b00000000 ;
			15'h00005765 : data <= 8'b00000000 ;
			15'h00005766 : data <= 8'b00000000 ;
			15'h00005767 : data <= 8'b00000000 ;
			15'h00005768 : data <= 8'b00000000 ;
			15'h00005769 : data <= 8'b00000000 ;
			15'h0000576A : data <= 8'b00000000 ;
			15'h0000576B : data <= 8'b00000000 ;
			15'h0000576C : data <= 8'b00000000 ;
			15'h0000576D : data <= 8'b00000000 ;
			15'h0000576E : data <= 8'b00000000 ;
			15'h0000576F : data <= 8'b00000000 ;
			15'h00005770 : data <= 8'b00000000 ;
			15'h00005771 : data <= 8'b00000000 ;
			15'h00005772 : data <= 8'b00000000 ;
			15'h00005773 : data <= 8'b00000000 ;
			15'h00005774 : data <= 8'b00000000 ;
			15'h00005775 : data <= 8'b00000000 ;
			15'h00005776 : data <= 8'b00000000 ;
			15'h00005777 : data <= 8'b00000000 ;
			15'h00005778 : data <= 8'b00000000 ;
			15'h00005779 : data <= 8'b00000000 ;
			15'h0000577A : data <= 8'b00000000 ;
			15'h0000577B : data <= 8'b00000000 ;
			15'h0000577C : data <= 8'b00000000 ;
			15'h0000577D : data <= 8'b00000000 ;
			15'h0000577E : data <= 8'b00000000 ;
			15'h0000577F : data <= 8'b00000000 ;
			15'h00005780 : data <= 8'b00000000 ;
			15'h00005781 : data <= 8'b00000000 ;
			15'h00005782 : data <= 8'b00000000 ;
			15'h00005783 : data <= 8'b00000000 ;
			15'h00005784 : data <= 8'b00000000 ;
			15'h00005785 : data <= 8'b00000000 ;
			15'h00005786 : data <= 8'b00000000 ;
			15'h00005787 : data <= 8'b00000000 ;
			15'h00005788 : data <= 8'b00000000 ;
			15'h00005789 : data <= 8'b00000000 ;
			15'h0000578A : data <= 8'b00000000 ;
			15'h0000578B : data <= 8'b00000000 ;
			15'h0000578C : data <= 8'b00000000 ;
			15'h0000578D : data <= 8'b00000000 ;
			15'h0000578E : data <= 8'b00000000 ;
			15'h0000578F : data <= 8'b00000000 ;
			15'h00005790 : data <= 8'b00000000 ;
			15'h00005791 : data <= 8'b00000000 ;
			15'h00005792 : data <= 8'b00000000 ;
			15'h00005793 : data <= 8'b00000000 ;
			15'h00005794 : data <= 8'b00000000 ;
			15'h00005795 : data <= 8'b00000000 ;
			15'h00005796 : data <= 8'b00000000 ;
			15'h00005797 : data <= 8'b00000000 ;
			15'h00005798 : data <= 8'b00000000 ;
			15'h00005799 : data <= 8'b00000000 ;
			15'h0000579A : data <= 8'b00000000 ;
			15'h0000579B : data <= 8'b00000000 ;
			15'h0000579C : data <= 8'b00000000 ;
			15'h0000579D : data <= 8'b00000000 ;
			15'h0000579E : data <= 8'b00000000 ;
			15'h0000579F : data <= 8'b00000000 ;
			15'h000057A0 : data <= 8'b00000000 ;
			15'h000057A1 : data <= 8'b00000000 ;
			15'h000057A2 : data <= 8'b00000000 ;
			15'h000057A3 : data <= 8'b00000000 ;
			15'h000057A4 : data <= 8'b00000000 ;
			15'h000057A5 : data <= 8'b00000000 ;
			15'h000057A6 : data <= 8'b00000000 ;
			15'h000057A7 : data <= 8'b00000000 ;
			15'h000057A8 : data <= 8'b00000000 ;
			15'h000057A9 : data <= 8'b00000000 ;
			15'h000057AA : data <= 8'b00000000 ;
			15'h000057AB : data <= 8'b00000000 ;
			15'h000057AC : data <= 8'b00000000 ;
			15'h000057AD : data <= 8'b00000000 ;
			15'h000057AE : data <= 8'b00000000 ;
			15'h000057AF : data <= 8'b00000000 ;
			15'h000057B0 : data <= 8'b00000000 ;
			15'h000057B1 : data <= 8'b00000000 ;
			15'h000057B2 : data <= 8'b00000000 ;
			15'h000057B3 : data <= 8'b00000000 ;
			15'h000057B4 : data <= 8'b00000000 ;
			15'h000057B5 : data <= 8'b00000000 ;
			15'h000057B6 : data <= 8'b00000000 ;
			15'h000057B7 : data <= 8'b00000000 ;
			15'h000057B8 : data <= 8'b00000000 ;
			15'h000057B9 : data <= 8'b00000000 ;
			15'h000057BA : data <= 8'b00000000 ;
			15'h000057BB : data <= 8'b00000000 ;
			15'h000057BC : data <= 8'b00000000 ;
			15'h000057BD : data <= 8'b00000000 ;
			15'h000057BE : data <= 8'b00000000 ;
			15'h000057BF : data <= 8'b00000000 ;
			15'h000057C0 : data <= 8'b00000000 ;
			15'h000057C1 : data <= 8'b00000000 ;
			15'h000057C2 : data <= 8'b00000000 ;
			15'h000057C3 : data <= 8'b00000000 ;
			15'h000057C4 : data <= 8'b00000000 ;
			15'h000057C5 : data <= 8'b00000000 ;
			15'h000057C6 : data <= 8'b00000000 ;
			15'h000057C7 : data <= 8'b00000000 ;
			15'h000057C8 : data <= 8'b00000000 ;
			15'h000057C9 : data <= 8'b00000000 ;
			15'h000057CA : data <= 8'b00000000 ;
			15'h000057CB : data <= 8'b00000000 ;
			15'h000057CC : data <= 8'b00000000 ;
			15'h000057CD : data <= 8'b00000000 ;
			15'h000057CE : data <= 8'b00000000 ;
			15'h000057CF : data <= 8'b00000000 ;
			15'h000057D0 : data <= 8'b00000000 ;
			15'h000057D1 : data <= 8'b00000000 ;
			15'h000057D2 : data <= 8'b00000000 ;
			15'h000057D3 : data <= 8'b00000000 ;
			15'h000057D4 : data <= 8'b00000000 ;
			15'h000057D5 : data <= 8'b00000000 ;
			15'h000057D6 : data <= 8'b00000000 ;
			15'h000057D7 : data <= 8'b00000000 ;
			15'h000057D8 : data <= 8'b00000000 ;
			15'h000057D9 : data <= 8'b00000000 ;
			15'h000057DA : data <= 8'b00000000 ;
			15'h000057DB : data <= 8'b00000000 ;
			15'h000057DC : data <= 8'b00000000 ;
			15'h000057DD : data <= 8'b00000000 ;
			15'h000057DE : data <= 8'b00000000 ;
			15'h000057DF : data <= 8'b00000000 ;
			15'h000057E0 : data <= 8'b00000000 ;
			15'h000057E1 : data <= 8'b00000000 ;
			15'h000057E2 : data <= 8'b00000000 ;
			15'h000057E3 : data <= 8'b00000000 ;
			15'h000057E4 : data <= 8'b00000000 ;
			15'h000057E5 : data <= 8'b00000000 ;
			15'h000057E6 : data <= 8'b00000000 ;
			15'h000057E7 : data <= 8'b00000000 ;
			15'h000057E8 : data <= 8'b00000000 ;
			15'h000057E9 : data <= 8'b00000000 ;
			15'h000057EA : data <= 8'b00000000 ;
			15'h000057EB : data <= 8'b00000000 ;
			15'h000057EC : data <= 8'b00000000 ;
			15'h000057ED : data <= 8'b00000000 ;
			15'h000057EE : data <= 8'b00000000 ;
			15'h000057EF : data <= 8'b00000000 ;
			15'h000057F0 : data <= 8'b00000000 ;
			15'h000057F1 : data <= 8'b00000000 ;
			15'h000057F2 : data <= 8'b00000000 ;
			15'h000057F3 : data <= 8'b00000000 ;
			15'h000057F4 : data <= 8'b00000000 ;
			15'h000057F5 : data <= 8'b00000000 ;
			15'h000057F6 : data <= 8'b00000000 ;
			15'h000057F7 : data <= 8'b00000000 ;
			15'h000057F8 : data <= 8'b00000000 ;
			15'h000057F9 : data <= 8'b00000000 ;
			15'h000057FA : data <= 8'b00000000 ;
			15'h000057FB : data <= 8'b00000000 ;
			15'h000057FC : data <= 8'b00000000 ;
			15'h000057FD : data <= 8'b00000000 ;
			15'h000057FE : data <= 8'b00000000 ;
			15'h000057FF : data <= 8'b00000000 ;
			15'h00005800 : data <= 8'b00000000 ;
			15'h00005801 : data <= 8'b00000000 ;
			15'h00005802 : data <= 8'b00000000 ;
			15'h00005803 : data <= 8'b00000000 ;
			15'h00005804 : data <= 8'b00000000 ;
			15'h00005805 : data <= 8'b00000000 ;
			15'h00005806 : data <= 8'b00000000 ;
			15'h00005807 : data <= 8'b00000000 ;
			15'h00005808 : data <= 8'b00000000 ;
			15'h00005809 : data <= 8'b00000000 ;
			15'h0000580A : data <= 8'b00000000 ;
			15'h0000580B : data <= 8'b00000000 ;
			15'h0000580C : data <= 8'b00000000 ;
			15'h0000580D : data <= 8'b00000000 ;
			15'h0000580E : data <= 8'b00000000 ;
			15'h0000580F : data <= 8'b00000000 ;
			15'h00005810 : data <= 8'b00000000 ;
			15'h00005811 : data <= 8'b00000000 ;
			15'h00005812 : data <= 8'b00000000 ;
			15'h00005813 : data <= 8'b00000000 ;
			15'h00005814 : data <= 8'b00000000 ;
			15'h00005815 : data <= 8'b00000000 ;
			15'h00005816 : data <= 8'b00000000 ;
			15'h00005817 : data <= 8'b00000000 ;
			15'h00005818 : data <= 8'b00000000 ;
			15'h00005819 : data <= 8'b00000000 ;
			15'h0000581A : data <= 8'b00000000 ;
			15'h0000581B : data <= 8'b00000000 ;
			15'h0000581C : data <= 8'b00000000 ;
			15'h0000581D : data <= 8'b00000000 ;
			15'h0000581E : data <= 8'b00000000 ;
			15'h0000581F : data <= 8'b00000000 ;
			15'h00005820 : data <= 8'b00000000 ;
			15'h00005821 : data <= 8'b00000000 ;
			15'h00005822 : data <= 8'b00000000 ;
			15'h00005823 : data <= 8'b00000000 ;
			15'h00005824 : data <= 8'b00000000 ;
			15'h00005825 : data <= 8'b00000000 ;
			15'h00005826 : data <= 8'b00000000 ;
			15'h00005827 : data <= 8'b00000000 ;
			15'h00005828 : data <= 8'b00000000 ;
			15'h00005829 : data <= 8'b00000000 ;
			15'h0000582A : data <= 8'b00000000 ;
			15'h0000582B : data <= 8'b00000000 ;
			15'h0000582C : data <= 8'b00000000 ;
			15'h0000582D : data <= 8'b00000000 ;
			15'h0000582E : data <= 8'b00000000 ;
			15'h0000582F : data <= 8'b00000000 ;
			15'h00005830 : data <= 8'b00000000 ;
			15'h00005831 : data <= 8'b00000000 ;
			15'h00005832 : data <= 8'b00000000 ;
			15'h00005833 : data <= 8'b00000000 ;
			15'h00005834 : data <= 8'b00000000 ;
			15'h00005835 : data <= 8'b00000000 ;
			15'h00005836 : data <= 8'b00000000 ;
			15'h00005837 : data <= 8'b00000000 ;
			15'h00005838 : data <= 8'b00000000 ;
			15'h00005839 : data <= 8'b00000000 ;
			15'h0000583A : data <= 8'b00000000 ;
			15'h0000583B : data <= 8'b00000000 ;
			15'h0000583C : data <= 8'b00000000 ;
			15'h0000583D : data <= 8'b00000000 ;
			15'h0000583E : data <= 8'b00000000 ;
			15'h0000583F : data <= 8'b00000000 ;
			15'h00005840 : data <= 8'b00000000 ;
			15'h00005841 : data <= 8'b00000000 ;
			15'h00005842 : data <= 8'b00000000 ;
			15'h00005843 : data <= 8'b00000000 ;
			15'h00005844 : data <= 8'b00000000 ;
			15'h00005845 : data <= 8'b00000000 ;
			15'h00005846 : data <= 8'b00000000 ;
			15'h00005847 : data <= 8'b00000000 ;
			15'h00005848 : data <= 8'b00000000 ;
			15'h00005849 : data <= 8'b00000000 ;
			15'h0000584A : data <= 8'b00000000 ;
			15'h0000584B : data <= 8'b00000000 ;
			15'h0000584C : data <= 8'b00000000 ;
			15'h0000584D : data <= 8'b00000000 ;
			15'h0000584E : data <= 8'b00000000 ;
			15'h0000584F : data <= 8'b00000000 ;
			15'h00005850 : data <= 8'b00000000 ;
			15'h00005851 : data <= 8'b00000000 ;
			15'h00005852 : data <= 8'b00000000 ;
			15'h00005853 : data <= 8'b00000000 ;
			15'h00005854 : data <= 8'b00000000 ;
			15'h00005855 : data <= 8'b00000000 ;
			15'h00005856 : data <= 8'b00000000 ;
			15'h00005857 : data <= 8'b00000000 ;
			15'h00005858 : data <= 8'b00000000 ;
			15'h00005859 : data <= 8'b00000000 ;
			15'h0000585A : data <= 8'b00000000 ;
			15'h0000585B : data <= 8'b00000000 ;
			15'h0000585C : data <= 8'b00000000 ;
			15'h0000585D : data <= 8'b00000000 ;
			15'h0000585E : data <= 8'b00000000 ;
			15'h0000585F : data <= 8'b00000000 ;
			15'h00005860 : data <= 8'b00000000 ;
			15'h00005861 : data <= 8'b00000000 ;
			15'h00005862 : data <= 8'b00000000 ;
			15'h00005863 : data <= 8'b00000000 ;
			15'h00005864 : data <= 8'b00000000 ;
			15'h00005865 : data <= 8'b00000000 ;
			15'h00005866 : data <= 8'b00000000 ;
			15'h00005867 : data <= 8'b00000000 ;
			15'h00005868 : data <= 8'b00000000 ;
			15'h00005869 : data <= 8'b00000000 ;
			15'h0000586A : data <= 8'b00000000 ;
			15'h0000586B : data <= 8'b00000000 ;
			15'h0000586C : data <= 8'b00000000 ;
			15'h0000586D : data <= 8'b00000000 ;
			15'h0000586E : data <= 8'b00000000 ;
			15'h0000586F : data <= 8'b00000000 ;
			15'h00005870 : data <= 8'b00000000 ;
			15'h00005871 : data <= 8'b00000000 ;
			15'h00005872 : data <= 8'b00000000 ;
			15'h00005873 : data <= 8'b00000000 ;
			15'h00005874 : data <= 8'b00000000 ;
			15'h00005875 : data <= 8'b00000000 ;
			15'h00005876 : data <= 8'b00000000 ;
			15'h00005877 : data <= 8'b00000000 ;
			15'h00005878 : data <= 8'b00000000 ;
			15'h00005879 : data <= 8'b00000000 ;
			15'h0000587A : data <= 8'b00000000 ;
			15'h0000587B : data <= 8'b00000000 ;
			15'h0000587C : data <= 8'b00000000 ;
			15'h0000587D : data <= 8'b00000000 ;
			15'h0000587E : data <= 8'b00000000 ;
			15'h0000587F : data <= 8'b00000000 ;
			15'h00005880 : data <= 8'b00000000 ;
			15'h00005881 : data <= 8'b00000000 ;
			15'h00005882 : data <= 8'b00000000 ;
			15'h00005883 : data <= 8'b00000000 ;
			15'h00005884 : data <= 8'b00000000 ;
			15'h00005885 : data <= 8'b00000000 ;
			15'h00005886 : data <= 8'b00000000 ;
			15'h00005887 : data <= 8'b00000000 ;
			15'h00005888 : data <= 8'b00000000 ;
			15'h00005889 : data <= 8'b00000000 ;
			15'h0000588A : data <= 8'b00000000 ;
			15'h0000588B : data <= 8'b00000000 ;
			15'h0000588C : data <= 8'b00000000 ;
			15'h0000588D : data <= 8'b00000000 ;
			15'h0000588E : data <= 8'b00000000 ;
			15'h0000588F : data <= 8'b00000000 ;
			15'h00005890 : data <= 8'b00000000 ;
			15'h00005891 : data <= 8'b00000000 ;
			15'h00005892 : data <= 8'b00000000 ;
			15'h00005893 : data <= 8'b00000000 ;
			15'h00005894 : data <= 8'b00000000 ;
			15'h00005895 : data <= 8'b00000000 ;
			15'h00005896 : data <= 8'b00000000 ;
			15'h00005897 : data <= 8'b00000000 ;
			15'h00005898 : data <= 8'b00000000 ;
			15'h00005899 : data <= 8'b00000000 ;
			15'h0000589A : data <= 8'b00000000 ;
			15'h0000589B : data <= 8'b00000000 ;
			15'h0000589C : data <= 8'b00000000 ;
			15'h0000589D : data <= 8'b00000000 ;
			15'h0000589E : data <= 8'b00000000 ;
			15'h0000589F : data <= 8'b00000000 ;
			15'h000058A0 : data <= 8'b00000000 ;
			15'h000058A1 : data <= 8'b00000000 ;
			15'h000058A2 : data <= 8'b00000000 ;
			15'h000058A3 : data <= 8'b00000000 ;
			15'h000058A4 : data <= 8'b00000000 ;
			15'h000058A5 : data <= 8'b00000000 ;
			15'h000058A6 : data <= 8'b00000000 ;
			15'h000058A7 : data <= 8'b00000000 ;
			15'h000058A8 : data <= 8'b00000000 ;
			15'h000058A9 : data <= 8'b00000000 ;
			15'h000058AA : data <= 8'b00000000 ;
			15'h000058AB : data <= 8'b00000000 ;
			15'h000058AC : data <= 8'b00000000 ;
			15'h000058AD : data <= 8'b00000000 ;
			15'h000058AE : data <= 8'b00000000 ;
			15'h000058AF : data <= 8'b00000000 ;
			15'h000058B0 : data <= 8'b00000000 ;
			15'h000058B1 : data <= 8'b00000000 ;
			15'h000058B2 : data <= 8'b00000000 ;
			15'h000058B3 : data <= 8'b00000000 ;
			15'h000058B4 : data <= 8'b00000000 ;
			15'h000058B5 : data <= 8'b00000000 ;
			15'h000058B6 : data <= 8'b00000000 ;
			15'h000058B7 : data <= 8'b00000000 ;
			15'h000058B8 : data <= 8'b00000000 ;
			15'h000058B9 : data <= 8'b00000000 ;
			15'h000058BA : data <= 8'b00000000 ;
			15'h000058BB : data <= 8'b00000000 ;
			15'h000058BC : data <= 8'b00000000 ;
			15'h000058BD : data <= 8'b00000000 ;
			15'h000058BE : data <= 8'b00000000 ;
			15'h000058BF : data <= 8'b00000000 ;
			15'h000058C0 : data <= 8'b00000000 ;
			15'h000058C1 : data <= 8'b00000000 ;
			15'h000058C2 : data <= 8'b00000000 ;
			15'h000058C3 : data <= 8'b00000000 ;
			15'h000058C4 : data <= 8'b00000000 ;
			15'h000058C5 : data <= 8'b00000000 ;
			15'h000058C6 : data <= 8'b00000000 ;
			15'h000058C7 : data <= 8'b00000000 ;
			15'h000058C8 : data <= 8'b00000000 ;
			15'h000058C9 : data <= 8'b00000000 ;
			15'h000058CA : data <= 8'b00000000 ;
			15'h000058CB : data <= 8'b00000000 ;
			15'h000058CC : data <= 8'b00000000 ;
			15'h000058CD : data <= 8'b00000000 ;
			15'h000058CE : data <= 8'b00000000 ;
			15'h000058CF : data <= 8'b00000000 ;
			15'h000058D0 : data <= 8'b00000000 ;
			15'h000058D1 : data <= 8'b00000000 ;
			15'h000058D2 : data <= 8'b00000000 ;
			15'h000058D3 : data <= 8'b00000000 ;
			15'h000058D4 : data <= 8'b00000000 ;
			15'h000058D5 : data <= 8'b00000000 ;
			15'h000058D6 : data <= 8'b00000000 ;
			15'h000058D7 : data <= 8'b00000000 ;
			15'h000058D8 : data <= 8'b00000000 ;
			15'h000058D9 : data <= 8'b00000000 ;
			15'h000058DA : data <= 8'b00000000 ;
			15'h000058DB : data <= 8'b00000000 ;
			15'h000058DC : data <= 8'b00000000 ;
			15'h000058DD : data <= 8'b00000000 ;
			15'h000058DE : data <= 8'b00000000 ;
			15'h000058DF : data <= 8'b00000000 ;
			15'h000058E0 : data <= 8'b00000000 ;
			15'h000058E1 : data <= 8'b00000000 ;
			15'h000058E2 : data <= 8'b00000000 ;
			15'h000058E3 : data <= 8'b00000000 ;
			15'h000058E4 : data <= 8'b00000000 ;
			15'h000058E5 : data <= 8'b00000000 ;
			15'h000058E6 : data <= 8'b00000000 ;
			15'h000058E7 : data <= 8'b00000000 ;
			15'h000058E8 : data <= 8'b00000000 ;
			15'h000058E9 : data <= 8'b00000000 ;
			15'h000058EA : data <= 8'b00000000 ;
			15'h000058EB : data <= 8'b00000000 ;
			15'h000058EC : data <= 8'b00000000 ;
			15'h000058ED : data <= 8'b00000000 ;
			15'h000058EE : data <= 8'b00000000 ;
			15'h000058EF : data <= 8'b00000000 ;
			15'h000058F0 : data <= 8'b00000000 ;
			15'h000058F1 : data <= 8'b00000000 ;
			15'h000058F2 : data <= 8'b00000000 ;
			15'h000058F3 : data <= 8'b00000000 ;
			15'h000058F4 : data <= 8'b00000000 ;
			15'h000058F5 : data <= 8'b00000000 ;
			15'h000058F6 : data <= 8'b00000000 ;
			15'h000058F7 : data <= 8'b00000000 ;
			15'h000058F8 : data <= 8'b00000000 ;
			15'h000058F9 : data <= 8'b00000000 ;
			15'h000058FA : data <= 8'b00000000 ;
			15'h000058FB : data <= 8'b00000000 ;
			15'h000058FC : data <= 8'b00000000 ;
			15'h000058FD : data <= 8'b00000000 ;
			15'h000058FE : data <= 8'b00000000 ;
			15'h000058FF : data <= 8'b00000000 ;
			15'h00005900 : data <= 8'b00000000 ;
			15'h00005901 : data <= 8'b00000000 ;
			15'h00005902 : data <= 8'b00000000 ;
			15'h00005903 : data <= 8'b00000000 ;
			15'h00005904 : data <= 8'b00000000 ;
			15'h00005905 : data <= 8'b00000000 ;
			15'h00005906 : data <= 8'b00000000 ;
			15'h00005907 : data <= 8'b00000000 ;
			15'h00005908 : data <= 8'b00000000 ;
			15'h00005909 : data <= 8'b00000000 ;
			15'h0000590A : data <= 8'b00000000 ;
			15'h0000590B : data <= 8'b00000000 ;
			15'h0000590C : data <= 8'b00000000 ;
			15'h0000590D : data <= 8'b00000000 ;
			15'h0000590E : data <= 8'b00000000 ;
			15'h0000590F : data <= 8'b00000000 ;
			15'h00005910 : data <= 8'b00000000 ;
			15'h00005911 : data <= 8'b00000000 ;
			15'h00005912 : data <= 8'b00000000 ;
			15'h00005913 : data <= 8'b00000000 ;
			15'h00005914 : data <= 8'b00000000 ;
			15'h00005915 : data <= 8'b00000000 ;
			15'h00005916 : data <= 8'b00000000 ;
			15'h00005917 : data <= 8'b00000000 ;
			15'h00005918 : data <= 8'b00000000 ;
			15'h00005919 : data <= 8'b00000000 ;
			15'h0000591A : data <= 8'b00000000 ;
			15'h0000591B : data <= 8'b00000000 ;
			15'h0000591C : data <= 8'b00000000 ;
			15'h0000591D : data <= 8'b00000000 ;
			15'h0000591E : data <= 8'b00000000 ;
			15'h0000591F : data <= 8'b00000000 ;
			15'h00005920 : data <= 8'b00000000 ;
			15'h00005921 : data <= 8'b00000000 ;
			15'h00005922 : data <= 8'b00000000 ;
			15'h00005923 : data <= 8'b00000000 ;
			15'h00005924 : data <= 8'b00000000 ;
			15'h00005925 : data <= 8'b00000000 ;
			15'h00005926 : data <= 8'b00000000 ;
			15'h00005927 : data <= 8'b00000000 ;
			15'h00005928 : data <= 8'b00000000 ;
			15'h00005929 : data <= 8'b00000000 ;
			15'h0000592A : data <= 8'b00000000 ;
			15'h0000592B : data <= 8'b00000000 ;
			15'h0000592C : data <= 8'b00000000 ;
			15'h0000592D : data <= 8'b00000000 ;
			15'h0000592E : data <= 8'b00000000 ;
			15'h0000592F : data <= 8'b00000000 ;
			15'h00005930 : data <= 8'b00000000 ;
			15'h00005931 : data <= 8'b00000000 ;
			15'h00005932 : data <= 8'b00000000 ;
			15'h00005933 : data <= 8'b00000000 ;
			15'h00005934 : data <= 8'b00000000 ;
			15'h00005935 : data <= 8'b00000000 ;
			15'h00005936 : data <= 8'b00000000 ;
			15'h00005937 : data <= 8'b00000000 ;
			15'h00005938 : data <= 8'b00000000 ;
			15'h00005939 : data <= 8'b00000000 ;
			15'h0000593A : data <= 8'b00000000 ;
			15'h0000593B : data <= 8'b00000000 ;
			15'h0000593C : data <= 8'b00000000 ;
			15'h0000593D : data <= 8'b00000000 ;
			15'h0000593E : data <= 8'b00000000 ;
			15'h0000593F : data <= 8'b00000000 ;
			15'h00005940 : data <= 8'b00000000 ;
			15'h00005941 : data <= 8'b00000000 ;
			15'h00005942 : data <= 8'b00000000 ;
			15'h00005943 : data <= 8'b00000000 ;
			15'h00005944 : data <= 8'b00000000 ;
			15'h00005945 : data <= 8'b00000000 ;
			15'h00005946 : data <= 8'b00000000 ;
			15'h00005947 : data <= 8'b00000000 ;
			15'h00005948 : data <= 8'b00000000 ;
			15'h00005949 : data <= 8'b00000000 ;
			15'h0000594A : data <= 8'b00000000 ;
			15'h0000594B : data <= 8'b00000000 ;
			15'h0000594C : data <= 8'b00000000 ;
			15'h0000594D : data <= 8'b00000000 ;
			15'h0000594E : data <= 8'b00000000 ;
			15'h0000594F : data <= 8'b00000000 ;
			15'h00005950 : data <= 8'b00000000 ;
			15'h00005951 : data <= 8'b00000000 ;
			15'h00005952 : data <= 8'b00000000 ;
			15'h00005953 : data <= 8'b00000000 ;
			15'h00005954 : data <= 8'b00000000 ;
			15'h00005955 : data <= 8'b00000000 ;
			15'h00005956 : data <= 8'b00000000 ;
			15'h00005957 : data <= 8'b00000000 ;
			15'h00005958 : data <= 8'b00000000 ;
			15'h00005959 : data <= 8'b00000000 ;
			15'h0000595A : data <= 8'b00000000 ;
			15'h0000595B : data <= 8'b00000000 ;
			15'h0000595C : data <= 8'b00000000 ;
			15'h0000595D : data <= 8'b00000000 ;
			15'h0000595E : data <= 8'b00000000 ;
			15'h0000595F : data <= 8'b00000000 ;
			15'h00005960 : data <= 8'b00000000 ;
			15'h00005961 : data <= 8'b00000000 ;
			15'h00005962 : data <= 8'b00000000 ;
			15'h00005963 : data <= 8'b00000000 ;
			15'h00005964 : data <= 8'b00000000 ;
			15'h00005965 : data <= 8'b00000000 ;
			15'h00005966 : data <= 8'b00000000 ;
			15'h00005967 : data <= 8'b00000000 ;
			15'h00005968 : data <= 8'b00000000 ;
			15'h00005969 : data <= 8'b00000000 ;
			15'h0000596A : data <= 8'b00000000 ;
			15'h0000596B : data <= 8'b00000000 ;
			15'h0000596C : data <= 8'b00000000 ;
			15'h0000596D : data <= 8'b00000000 ;
			15'h0000596E : data <= 8'b00000000 ;
			15'h0000596F : data <= 8'b00000000 ;
			15'h00005970 : data <= 8'b00000000 ;
			15'h00005971 : data <= 8'b00000000 ;
			15'h00005972 : data <= 8'b00000000 ;
			15'h00005973 : data <= 8'b00000000 ;
			15'h00005974 : data <= 8'b00000000 ;
			15'h00005975 : data <= 8'b00000000 ;
			15'h00005976 : data <= 8'b00000000 ;
			15'h00005977 : data <= 8'b00000000 ;
			15'h00005978 : data <= 8'b00000000 ;
			15'h00005979 : data <= 8'b00000000 ;
			15'h0000597A : data <= 8'b00000000 ;
			15'h0000597B : data <= 8'b00000000 ;
			15'h0000597C : data <= 8'b00000000 ;
			15'h0000597D : data <= 8'b00000000 ;
			15'h0000597E : data <= 8'b00000000 ;
			15'h0000597F : data <= 8'b00000000 ;
			15'h00005980 : data <= 8'b00000000 ;
			15'h00005981 : data <= 8'b00000000 ;
			15'h00005982 : data <= 8'b00000000 ;
			15'h00005983 : data <= 8'b00000000 ;
			15'h00005984 : data <= 8'b00000000 ;
			15'h00005985 : data <= 8'b00000000 ;
			15'h00005986 : data <= 8'b00000000 ;
			15'h00005987 : data <= 8'b00000000 ;
			15'h00005988 : data <= 8'b00000000 ;
			15'h00005989 : data <= 8'b00000000 ;
			15'h0000598A : data <= 8'b00000000 ;
			15'h0000598B : data <= 8'b00000000 ;
			15'h0000598C : data <= 8'b00000000 ;
			15'h0000598D : data <= 8'b00000000 ;
			15'h0000598E : data <= 8'b00000000 ;
			15'h0000598F : data <= 8'b00000000 ;
			15'h00005990 : data <= 8'b00000000 ;
			15'h00005991 : data <= 8'b00000000 ;
			15'h00005992 : data <= 8'b00000000 ;
			15'h00005993 : data <= 8'b00000000 ;
			15'h00005994 : data <= 8'b00000000 ;
			15'h00005995 : data <= 8'b00000000 ;
			15'h00005996 : data <= 8'b00000000 ;
			15'h00005997 : data <= 8'b00000000 ;
			15'h00005998 : data <= 8'b00000000 ;
			15'h00005999 : data <= 8'b00000000 ;
			15'h0000599A : data <= 8'b00000000 ;
			15'h0000599B : data <= 8'b00000000 ;
			15'h0000599C : data <= 8'b00000000 ;
			15'h0000599D : data <= 8'b00000000 ;
			15'h0000599E : data <= 8'b00000000 ;
			15'h0000599F : data <= 8'b00000000 ;
			15'h000059A0 : data <= 8'b00000000 ;
			15'h000059A1 : data <= 8'b00000000 ;
			15'h000059A2 : data <= 8'b00000000 ;
			15'h000059A3 : data <= 8'b00000000 ;
			15'h000059A4 : data <= 8'b00000000 ;
			15'h000059A5 : data <= 8'b00000000 ;
			15'h000059A6 : data <= 8'b00000000 ;
			15'h000059A7 : data <= 8'b00000000 ;
			15'h000059A8 : data <= 8'b00000000 ;
			15'h000059A9 : data <= 8'b00000000 ;
			15'h000059AA : data <= 8'b00000000 ;
			15'h000059AB : data <= 8'b00000000 ;
			15'h000059AC : data <= 8'b00000000 ;
			15'h000059AD : data <= 8'b00000000 ;
			15'h000059AE : data <= 8'b00000000 ;
			15'h000059AF : data <= 8'b00000000 ;
			15'h000059B0 : data <= 8'b00000000 ;
			15'h000059B1 : data <= 8'b00000000 ;
			15'h000059B2 : data <= 8'b00000000 ;
			15'h000059B3 : data <= 8'b00000000 ;
			15'h000059B4 : data <= 8'b00000000 ;
			15'h000059B5 : data <= 8'b00000000 ;
			15'h000059B6 : data <= 8'b00000000 ;
			15'h000059B7 : data <= 8'b00000000 ;
			15'h000059B8 : data <= 8'b00000000 ;
			15'h000059B9 : data <= 8'b00000000 ;
			15'h000059BA : data <= 8'b00000000 ;
			15'h000059BB : data <= 8'b00000000 ;
			15'h000059BC : data <= 8'b00000000 ;
			15'h000059BD : data <= 8'b00000000 ;
			15'h000059BE : data <= 8'b00000000 ;
			15'h000059BF : data <= 8'b00000000 ;
			15'h000059C0 : data <= 8'b00000000 ;
			15'h000059C1 : data <= 8'b00000000 ;
			15'h000059C2 : data <= 8'b00000000 ;
			15'h000059C3 : data <= 8'b00000000 ;
			15'h000059C4 : data <= 8'b00000000 ;
			15'h000059C5 : data <= 8'b00000000 ;
			15'h000059C6 : data <= 8'b00000000 ;
			15'h000059C7 : data <= 8'b00000000 ;
			15'h000059C8 : data <= 8'b00000000 ;
			15'h000059C9 : data <= 8'b00000000 ;
			15'h000059CA : data <= 8'b00000000 ;
			15'h000059CB : data <= 8'b00000000 ;
			15'h000059CC : data <= 8'b00000000 ;
			15'h000059CD : data <= 8'b00000000 ;
			15'h000059CE : data <= 8'b00000000 ;
			15'h000059CF : data <= 8'b00000000 ;
			15'h000059D0 : data <= 8'b00000000 ;
			15'h000059D1 : data <= 8'b00000000 ;
			15'h000059D2 : data <= 8'b00000000 ;
			15'h000059D3 : data <= 8'b00000000 ;
			15'h000059D4 : data <= 8'b00000000 ;
			15'h000059D5 : data <= 8'b00000000 ;
			15'h000059D6 : data <= 8'b00000000 ;
			15'h000059D7 : data <= 8'b00000000 ;
			15'h000059D8 : data <= 8'b00000000 ;
			15'h000059D9 : data <= 8'b00000000 ;
			15'h000059DA : data <= 8'b00000000 ;
			15'h000059DB : data <= 8'b00000000 ;
			15'h000059DC : data <= 8'b00000000 ;
			15'h000059DD : data <= 8'b00000000 ;
			15'h000059DE : data <= 8'b00000000 ;
			15'h000059DF : data <= 8'b00000000 ;
			15'h000059E0 : data <= 8'b00000000 ;
			15'h000059E1 : data <= 8'b00000000 ;
			15'h000059E2 : data <= 8'b00000000 ;
			15'h000059E3 : data <= 8'b00000000 ;
			15'h000059E4 : data <= 8'b00000000 ;
			15'h000059E5 : data <= 8'b00000000 ;
			15'h000059E6 : data <= 8'b00000000 ;
			15'h000059E7 : data <= 8'b00000000 ;
			15'h000059E8 : data <= 8'b00000000 ;
			15'h000059E9 : data <= 8'b00000000 ;
			15'h000059EA : data <= 8'b00000000 ;
			15'h000059EB : data <= 8'b00000000 ;
			15'h000059EC : data <= 8'b00000000 ;
			15'h000059ED : data <= 8'b00000000 ;
			15'h000059EE : data <= 8'b00000000 ;
			15'h000059EF : data <= 8'b00000000 ;
			15'h000059F0 : data <= 8'b00000000 ;
			15'h000059F1 : data <= 8'b00000000 ;
			15'h000059F2 : data <= 8'b00000000 ;
			15'h000059F3 : data <= 8'b00000000 ;
			15'h000059F4 : data <= 8'b00000000 ;
			15'h000059F5 : data <= 8'b00000000 ;
			15'h000059F6 : data <= 8'b00000000 ;
			15'h000059F7 : data <= 8'b00000000 ;
			15'h000059F8 : data <= 8'b00000000 ;
			15'h000059F9 : data <= 8'b00000000 ;
			15'h000059FA : data <= 8'b00000000 ;
			15'h000059FB : data <= 8'b00000000 ;
			15'h000059FC : data <= 8'b00000000 ;
			15'h000059FD : data <= 8'b00000000 ;
			15'h000059FE : data <= 8'b00000000 ;
			15'h000059FF : data <= 8'b00000000 ;
			15'h00005A00 : data <= 8'b00000000 ;
			15'h00005A01 : data <= 8'b00000000 ;
			15'h00005A02 : data <= 8'b00000000 ;
			15'h00005A03 : data <= 8'b00000000 ;
			15'h00005A04 : data <= 8'b00000000 ;
			15'h00005A05 : data <= 8'b00000000 ;
			15'h00005A06 : data <= 8'b00000000 ;
			15'h00005A07 : data <= 8'b00000000 ;
			15'h00005A08 : data <= 8'b00000000 ;
			15'h00005A09 : data <= 8'b00000000 ;
			15'h00005A0A : data <= 8'b00000000 ;
			15'h00005A0B : data <= 8'b00000000 ;
			15'h00005A0C : data <= 8'b00000000 ;
			15'h00005A0D : data <= 8'b00000000 ;
			15'h00005A0E : data <= 8'b00000000 ;
			15'h00005A0F : data <= 8'b00000000 ;
			15'h00005A10 : data <= 8'b00000000 ;
			15'h00005A11 : data <= 8'b00000000 ;
			15'h00005A12 : data <= 8'b00000000 ;
			15'h00005A13 : data <= 8'b00000000 ;
			15'h00005A14 : data <= 8'b00000000 ;
			15'h00005A15 : data <= 8'b00000000 ;
			15'h00005A16 : data <= 8'b00000000 ;
			15'h00005A17 : data <= 8'b00000000 ;
			15'h00005A18 : data <= 8'b00000000 ;
			15'h00005A19 : data <= 8'b00000000 ;
			15'h00005A1A : data <= 8'b00000000 ;
			15'h00005A1B : data <= 8'b00000000 ;
			15'h00005A1C : data <= 8'b00000000 ;
			15'h00005A1D : data <= 8'b00000000 ;
			15'h00005A1E : data <= 8'b00000000 ;
			15'h00005A1F : data <= 8'b00000000 ;
			15'h00005A20 : data <= 8'b00000000 ;
			15'h00005A21 : data <= 8'b00000000 ;
			15'h00005A22 : data <= 8'b00000000 ;
			15'h00005A23 : data <= 8'b00000000 ;
			15'h00005A24 : data <= 8'b00000000 ;
			15'h00005A25 : data <= 8'b00000000 ;
			15'h00005A26 : data <= 8'b00000000 ;
			15'h00005A27 : data <= 8'b00000000 ;
			15'h00005A28 : data <= 8'b00000000 ;
			15'h00005A29 : data <= 8'b00000000 ;
			15'h00005A2A : data <= 8'b00000000 ;
			15'h00005A2B : data <= 8'b00000000 ;
			15'h00005A2C : data <= 8'b00000000 ;
			15'h00005A2D : data <= 8'b00000000 ;
			15'h00005A2E : data <= 8'b00000000 ;
			15'h00005A2F : data <= 8'b00000000 ;
			15'h00005A30 : data <= 8'b00000000 ;
			15'h00005A31 : data <= 8'b00000000 ;
			15'h00005A32 : data <= 8'b00000000 ;
			15'h00005A33 : data <= 8'b00000000 ;
			15'h00005A34 : data <= 8'b00000000 ;
			15'h00005A35 : data <= 8'b00000000 ;
			15'h00005A36 : data <= 8'b00000000 ;
			15'h00005A37 : data <= 8'b00000000 ;
			15'h00005A38 : data <= 8'b00000000 ;
			15'h00005A39 : data <= 8'b00000000 ;
			15'h00005A3A : data <= 8'b00000000 ;
			15'h00005A3B : data <= 8'b00000000 ;
			15'h00005A3C : data <= 8'b00000000 ;
			15'h00005A3D : data <= 8'b00000000 ;
			15'h00005A3E : data <= 8'b00000000 ;
			15'h00005A3F : data <= 8'b00000000 ;
			15'h00005A40 : data <= 8'b00000000 ;
			15'h00005A41 : data <= 8'b00000000 ;
			15'h00005A42 : data <= 8'b00000000 ;
			15'h00005A43 : data <= 8'b00000000 ;
			15'h00005A44 : data <= 8'b00000000 ;
			15'h00005A45 : data <= 8'b00000000 ;
			15'h00005A46 : data <= 8'b00000000 ;
			15'h00005A47 : data <= 8'b00000000 ;
			15'h00005A48 : data <= 8'b00000000 ;
			15'h00005A49 : data <= 8'b00000000 ;
			15'h00005A4A : data <= 8'b00000000 ;
			15'h00005A4B : data <= 8'b00000000 ;
			15'h00005A4C : data <= 8'b00000000 ;
			15'h00005A4D : data <= 8'b00000000 ;
			15'h00005A4E : data <= 8'b00000000 ;
			15'h00005A4F : data <= 8'b00000000 ;
			15'h00005A50 : data <= 8'b00000000 ;
			15'h00005A51 : data <= 8'b00000000 ;
			15'h00005A52 : data <= 8'b00000000 ;
			15'h00005A53 : data <= 8'b00000000 ;
			15'h00005A54 : data <= 8'b00000000 ;
			15'h00005A55 : data <= 8'b00000000 ;
			15'h00005A56 : data <= 8'b00000000 ;
			15'h00005A57 : data <= 8'b00000000 ;
			15'h00005A58 : data <= 8'b00000000 ;
			15'h00005A59 : data <= 8'b00000000 ;
			15'h00005A5A : data <= 8'b00000000 ;
			15'h00005A5B : data <= 8'b00000000 ;
			15'h00005A5C : data <= 8'b00000000 ;
			15'h00005A5D : data <= 8'b00000000 ;
			15'h00005A5E : data <= 8'b00000000 ;
			15'h00005A5F : data <= 8'b00000000 ;
			15'h00005A60 : data <= 8'b00000000 ;
			15'h00005A61 : data <= 8'b00000000 ;
			15'h00005A62 : data <= 8'b00000000 ;
			15'h00005A63 : data <= 8'b00000000 ;
			15'h00005A64 : data <= 8'b00000000 ;
			15'h00005A65 : data <= 8'b00000000 ;
			15'h00005A66 : data <= 8'b00000000 ;
			15'h00005A67 : data <= 8'b00000000 ;
			15'h00005A68 : data <= 8'b00000000 ;
			15'h00005A69 : data <= 8'b00000000 ;
			15'h00005A6A : data <= 8'b00000000 ;
			15'h00005A6B : data <= 8'b00000000 ;
			15'h00005A6C : data <= 8'b00000000 ;
			15'h00005A6D : data <= 8'b00000000 ;
			15'h00005A6E : data <= 8'b00000000 ;
			15'h00005A6F : data <= 8'b00000000 ;
			15'h00005A70 : data <= 8'b00000000 ;
			15'h00005A71 : data <= 8'b00000000 ;
			15'h00005A72 : data <= 8'b00000000 ;
			15'h00005A73 : data <= 8'b00000000 ;
			15'h00005A74 : data <= 8'b00000000 ;
			15'h00005A75 : data <= 8'b00000000 ;
			15'h00005A76 : data <= 8'b00000000 ;
			15'h00005A77 : data <= 8'b00000000 ;
			15'h00005A78 : data <= 8'b00000000 ;
			15'h00005A79 : data <= 8'b00000000 ;
			15'h00005A7A : data <= 8'b00000000 ;
			15'h00005A7B : data <= 8'b00000000 ;
			15'h00005A7C : data <= 8'b00000000 ;
			15'h00005A7D : data <= 8'b00000000 ;
			15'h00005A7E : data <= 8'b00000000 ;
			15'h00005A7F : data <= 8'b00000000 ;
			15'h00005A80 : data <= 8'b00000000 ;
			15'h00005A81 : data <= 8'b00000000 ;
			15'h00005A82 : data <= 8'b00000000 ;
			15'h00005A83 : data <= 8'b00000000 ;
			15'h00005A84 : data <= 8'b00000000 ;
			15'h00005A85 : data <= 8'b00000000 ;
			15'h00005A86 : data <= 8'b00000000 ;
			15'h00005A87 : data <= 8'b00000000 ;
			15'h00005A88 : data <= 8'b00000000 ;
			15'h00005A89 : data <= 8'b00000000 ;
			15'h00005A8A : data <= 8'b00000000 ;
			15'h00005A8B : data <= 8'b00000000 ;
			15'h00005A8C : data <= 8'b00000000 ;
			15'h00005A8D : data <= 8'b00000000 ;
			15'h00005A8E : data <= 8'b00000000 ;
			15'h00005A8F : data <= 8'b00000000 ;
			15'h00005A90 : data <= 8'b00000000 ;
			15'h00005A91 : data <= 8'b00000000 ;
			15'h00005A92 : data <= 8'b00000000 ;
			15'h00005A93 : data <= 8'b00000000 ;
			15'h00005A94 : data <= 8'b00000000 ;
			15'h00005A95 : data <= 8'b00000000 ;
			15'h00005A96 : data <= 8'b00000000 ;
			15'h00005A97 : data <= 8'b00000000 ;
			15'h00005A98 : data <= 8'b00000000 ;
			15'h00005A99 : data <= 8'b00000000 ;
			15'h00005A9A : data <= 8'b00000000 ;
			15'h00005A9B : data <= 8'b00000000 ;
			15'h00005A9C : data <= 8'b00000000 ;
			15'h00005A9D : data <= 8'b00000000 ;
			15'h00005A9E : data <= 8'b00000000 ;
			15'h00005A9F : data <= 8'b00000000 ;
			15'h00005AA0 : data <= 8'b00000000 ;
			15'h00005AA1 : data <= 8'b00000000 ;
			15'h00005AA2 : data <= 8'b00000000 ;
			15'h00005AA3 : data <= 8'b00000000 ;
			15'h00005AA4 : data <= 8'b00000000 ;
			15'h00005AA5 : data <= 8'b00000000 ;
			15'h00005AA6 : data <= 8'b00000000 ;
			15'h00005AA7 : data <= 8'b00000000 ;
			15'h00005AA8 : data <= 8'b00000000 ;
			15'h00005AA9 : data <= 8'b00000000 ;
			15'h00005AAA : data <= 8'b00000000 ;
			15'h00005AAB : data <= 8'b00000000 ;
			15'h00005AAC : data <= 8'b00000000 ;
			15'h00005AAD : data <= 8'b00000000 ;
			15'h00005AAE : data <= 8'b00000000 ;
			15'h00005AAF : data <= 8'b00000000 ;
			15'h00005AB0 : data <= 8'b00000000 ;
			15'h00005AB1 : data <= 8'b00000000 ;
			15'h00005AB2 : data <= 8'b00000000 ;
			15'h00005AB3 : data <= 8'b00000000 ;
			15'h00005AB4 : data <= 8'b00000000 ;
			15'h00005AB5 : data <= 8'b00000000 ;
			15'h00005AB6 : data <= 8'b00000000 ;
			15'h00005AB7 : data <= 8'b00000000 ;
			15'h00005AB8 : data <= 8'b00000000 ;
			15'h00005AB9 : data <= 8'b00000000 ;
			15'h00005ABA : data <= 8'b00000000 ;
			15'h00005ABB : data <= 8'b00000000 ;
			15'h00005ABC : data <= 8'b00000000 ;
			15'h00005ABD : data <= 8'b00000000 ;
			15'h00005ABE : data <= 8'b00000000 ;
			15'h00005ABF : data <= 8'b00000000 ;
			15'h00005AC0 : data <= 8'b00000000 ;
			15'h00005AC1 : data <= 8'b00000000 ;
			15'h00005AC2 : data <= 8'b00000000 ;
			15'h00005AC3 : data <= 8'b00000000 ;
			15'h00005AC4 : data <= 8'b00000000 ;
			15'h00005AC5 : data <= 8'b00000000 ;
			15'h00005AC6 : data <= 8'b00000000 ;
			15'h00005AC7 : data <= 8'b00000000 ;
			15'h00005AC8 : data <= 8'b00000000 ;
			15'h00005AC9 : data <= 8'b00000000 ;
			15'h00005ACA : data <= 8'b00000000 ;
			15'h00005ACB : data <= 8'b00000000 ;
			15'h00005ACC : data <= 8'b00000000 ;
			15'h00005ACD : data <= 8'b00000000 ;
			15'h00005ACE : data <= 8'b00000000 ;
			15'h00005ACF : data <= 8'b00000000 ;
			15'h00005AD0 : data <= 8'b00000000 ;
			15'h00005AD1 : data <= 8'b00000000 ;
			15'h00005AD2 : data <= 8'b00000000 ;
			15'h00005AD3 : data <= 8'b00000000 ;
			15'h00005AD4 : data <= 8'b00000000 ;
			15'h00005AD5 : data <= 8'b00000000 ;
			15'h00005AD6 : data <= 8'b00000000 ;
			15'h00005AD7 : data <= 8'b00000000 ;
			15'h00005AD8 : data <= 8'b00000000 ;
			15'h00005AD9 : data <= 8'b00000000 ;
			15'h00005ADA : data <= 8'b00000000 ;
			15'h00005ADB : data <= 8'b00000000 ;
			15'h00005ADC : data <= 8'b00000000 ;
			15'h00005ADD : data <= 8'b00000000 ;
			15'h00005ADE : data <= 8'b00000000 ;
			15'h00005ADF : data <= 8'b00000000 ;
			15'h00005AE0 : data <= 8'b00000000 ;
			15'h00005AE1 : data <= 8'b00000000 ;
			15'h00005AE2 : data <= 8'b00000000 ;
			15'h00005AE3 : data <= 8'b00000000 ;
			15'h00005AE4 : data <= 8'b00000000 ;
			15'h00005AE5 : data <= 8'b00000000 ;
			15'h00005AE6 : data <= 8'b00000000 ;
			15'h00005AE7 : data <= 8'b00000000 ;
			15'h00005AE8 : data <= 8'b00000000 ;
			15'h00005AE9 : data <= 8'b00000000 ;
			15'h00005AEA : data <= 8'b00000000 ;
			15'h00005AEB : data <= 8'b00000000 ;
			15'h00005AEC : data <= 8'b00000000 ;
			15'h00005AED : data <= 8'b00000000 ;
			15'h00005AEE : data <= 8'b00000000 ;
			15'h00005AEF : data <= 8'b00000000 ;
			15'h00005AF0 : data <= 8'b00000000 ;
			15'h00005AF1 : data <= 8'b00000000 ;
			15'h00005AF2 : data <= 8'b00000000 ;
			15'h00005AF3 : data <= 8'b00000000 ;
			15'h00005AF4 : data <= 8'b00000000 ;
			15'h00005AF5 : data <= 8'b00000000 ;
			15'h00005AF6 : data <= 8'b00000000 ;
			15'h00005AF7 : data <= 8'b00000000 ;
			15'h00005AF8 : data <= 8'b00000000 ;
			15'h00005AF9 : data <= 8'b00000000 ;
			15'h00005AFA : data <= 8'b00000000 ;
			15'h00005AFB : data <= 8'b00000000 ;
			15'h00005AFC : data <= 8'b00000000 ;
			15'h00005AFD : data <= 8'b00000000 ;
			15'h00005AFE : data <= 8'b00000000 ;
			15'h00005AFF : data <= 8'b00000000 ;
			15'h00005B00 : data <= 8'b00000000 ;
			15'h00005B01 : data <= 8'b00000000 ;
			15'h00005B02 : data <= 8'b00000000 ;
			15'h00005B03 : data <= 8'b00000000 ;
			15'h00005B04 : data <= 8'b00000000 ;
			15'h00005B05 : data <= 8'b00000000 ;
			15'h00005B06 : data <= 8'b00000000 ;
			15'h00005B07 : data <= 8'b00000000 ;
			15'h00005B08 : data <= 8'b00000000 ;
			15'h00005B09 : data <= 8'b00000000 ;
			15'h00005B0A : data <= 8'b00000000 ;
			15'h00005B0B : data <= 8'b00000000 ;
			15'h00005B0C : data <= 8'b00000000 ;
			15'h00005B0D : data <= 8'b00000000 ;
			15'h00005B0E : data <= 8'b00000000 ;
			15'h00005B0F : data <= 8'b00000000 ;
			15'h00005B10 : data <= 8'b00000000 ;
			15'h00005B11 : data <= 8'b00000000 ;
			15'h00005B12 : data <= 8'b00000000 ;
			15'h00005B13 : data <= 8'b00000000 ;
			15'h00005B14 : data <= 8'b00000000 ;
			15'h00005B15 : data <= 8'b00000000 ;
			15'h00005B16 : data <= 8'b00000000 ;
			15'h00005B17 : data <= 8'b00000000 ;
			15'h00005B18 : data <= 8'b00000000 ;
			15'h00005B19 : data <= 8'b00000000 ;
			15'h00005B1A : data <= 8'b00000000 ;
			15'h00005B1B : data <= 8'b00000000 ;
			15'h00005B1C : data <= 8'b00000000 ;
			15'h00005B1D : data <= 8'b00000000 ;
			15'h00005B1E : data <= 8'b00000000 ;
			15'h00005B1F : data <= 8'b00000000 ;
			15'h00005B20 : data <= 8'b00000000 ;
			15'h00005B21 : data <= 8'b00000000 ;
			15'h00005B22 : data <= 8'b00000000 ;
			15'h00005B23 : data <= 8'b00000000 ;
			15'h00005B24 : data <= 8'b00000000 ;
			15'h00005B25 : data <= 8'b00000000 ;
			15'h00005B26 : data <= 8'b00000000 ;
			15'h00005B27 : data <= 8'b00000000 ;
			15'h00005B28 : data <= 8'b00000000 ;
			15'h00005B29 : data <= 8'b00000000 ;
			15'h00005B2A : data <= 8'b00000000 ;
			15'h00005B2B : data <= 8'b00000000 ;
			15'h00005B2C : data <= 8'b00000000 ;
			15'h00005B2D : data <= 8'b00000000 ;
			15'h00005B2E : data <= 8'b00000000 ;
			15'h00005B2F : data <= 8'b00000000 ;
			15'h00005B30 : data <= 8'b00000000 ;
			15'h00005B31 : data <= 8'b00000000 ;
			15'h00005B32 : data <= 8'b00000000 ;
			15'h00005B33 : data <= 8'b00000000 ;
			15'h00005B34 : data <= 8'b00000000 ;
			15'h00005B35 : data <= 8'b00000000 ;
			15'h00005B36 : data <= 8'b00000000 ;
			15'h00005B37 : data <= 8'b00000000 ;
			15'h00005B38 : data <= 8'b00000000 ;
			15'h00005B39 : data <= 8'b00000000 ;
			15'h00005B3A : data <= 8'b00000000 ;
			15'h00005B3B : data <= 8'b00000000 ;
			15'h00005B3C : data <= 8'b00000000 ;
			15'h00005B3D : data <= 8'b00000000 ;
			15'h00005B3E : data <= 8'b00000000 ;
			15'h00005B3F : data <= 8'b00000000 ;
			15'h00005B40 : data <= 8'b00000000 ;
			15'h00005B41 : data <= 8'b00000000 ;
			15'h00005B42 : data <= 8'b00000000 ;
			15'h00005B43 : data <= 8'b00000000 ;
			15'h00005B44 : data <= 8'b00000000 ;
			15'h00005B45 : data <= 8'b00000000 ;
			15'h00005B46 : data <= 8'b00000000 ;
			15'h00005B47 : data <= 8'b00000000 ;
			15'h00005B48 : data <= 8'b00000000 ;
			15'h00005B49 : data <= 8'b00000000 ;
			15'h00005B4A : data <= 8'b00000000 ;
			15'h00005B4B : data <= 8'b00000000 ;
			15'h00005B4C : data <= 8'b00000000 ;
			15'h00005B4D : data <= 8'b00000000 ;
			15'h00005B4E : data <= 8'b00000000 ;
			15'h00005B4F : data <= 8'b00000000 ;
			15'h00005B50 : data <= 8'b00000000 ;
			15'h00005B51 : data <= 8'b00000000 ;
			15'h00005B52 : data <= 8'b00000000 ;
			15'h00005B53 : data <= 8'b00000000 ;
			15'h00005B54 : data <= 8'b00000000 ;
			15'h00005B55 : data <= 8'b00000000 ;
			15'h00005B56 : data <= 8'b00000000 ;
			15'h00005B57 : data <= 8'b00000000 ;
			15'h00005B58 : data <= 8'b00000000 ;
			15'h00005B59 : data <= 8'b00000000 ;
			15'h00005B5A : data <= 8'b00000000 ;
			15'h00005B5B : data <= 8'b00000000 ;
			15'h00005B5C : data <= 8'b00000000 ;
			15'h00005B5D : data <= 8'b00000000 ;
			15'h00005B5E : data <= 8'b00000000 ;
			15'h00005B5F : data <= 8'b00000000 ;
			15'h00005B60 : data <= 8'b00000000 ;
			15'h00005B61 : data <= 8'b00000000 ;
			15'h00005B62 : data <= 8'b00000000 ;
			15'h00005B63 : data <= 8'b00000000 ;
			15'h00005B64 : data <= 8'b00000000 ;
			15'h00005B65 : data <= 8'b00000000 ;
			15'h00005B66 : data <= 8'b00000000 ;
			15'h00005B67 : data <= 8'b00000000 ;
			15'h00005B68 : data <= 8'b00000000 ;
			15'h00005B69 : data <= 8'b00000000 ;
			15'h00005B6A : data <= 8'b00000000 ;
			15'h00005B6B : data <= 8'b00000000 ;
			15'h00005B6C : data <= 8'b00000000 ;
			15'h00005B6D : data <= 8'b00000000 ;
			15'h00005B6E : data <= 8'b00000000 ;
			15'h00005B6F : data <= 8'b00000000 ;
			15'h00005B70 : data <= 8'b00000000 ;
			15'h00005B71 : data <= 8'b00000000 ;
			15'h00005B72 : data <= 8'b00000000 ;
			15'h00005B73 : data <= 8'b00000000 ;
			15'h00005B74 : data <= 8'b00000000 ;
			15'h00005B75 : data <= 8'b00000000 ;
			15'h00005B76 : data <= 8'b00000000 ;
			15'h00005B77 : data <= 8'b00000000 ;
			15'h00005B78 : data <= 8'b00000000 ;
			15'h00005B79 : data <= 8'b00000000 ;
			15'h00005B7A : data <= 8'b00000000 ;
			15'h00005B7B : data <= 8'b00000000 ;
			15'h00005B7C : data <= 8'b00000000 ;
			15'h00005B7D : data <= 8'b00000000 ;
			15'h00005B7E : data <= 8'b00000000 ;
			15'h00005B7F : data <= 8'b00000000 ;
			15'h00005B80 : data <= 8'b00000000 ;
			15'h00005B81 : data <= 8'b00000000 ;
			15'h00005B82 : data <= 8'b00000000 ;
			15'h00005B83 : data <= 8'b00000000 ;
			15'h00005B84 : data <= 8'b00000000 ;
			15'h00005B85 : data <= 8'b00000000 ;
			15'h00005B86 : data <= 8'b00000000 ;
			15'h00005B87 : data <= 8'b00000000 ;
			15'h00005B88 : data <= 8'b00000000 ;
			15'h00005B89 : data <= 8'b00000000 ;
			15'h00005B8A : data <= 8'b00000000 ;
			15'h00005B8B : data <= 8'b00000000 ;
			15'h00005B8C : data <= 8'b00000000 ;
			15'h00005B8D : data <= 8'b00000000 ;
			15'h00005B8E : data <= 8'b00000000 ;
			15'h00005B8F : data <= 8'b00000000 ;
			15'h00005B90 : data <= 8'b00000000 ;
			15'h00005B91 : data <= 8'b00000000 ;
			15'h00005B92 : data <= 8'b00000000 ;
			15'h00005B93 : data <= 8'b00000000 ;
			15'h00005B94 : data <= 8'b00000000 ;
			15'h00005B95 : data <= 8'b00000000 ;
			15'h00005B96 : data <= 8'b00000000 ;
			15'h00005B97 : data <= 8'b00000000 ;
			15'h00005B98 : data <= 8'b00000000 ;
			15'h00005B99 : data <= 8'b00000000 ;
			15'h00005B9A : data <= 8'b00000000 ;
			15'h00005B9B : data <= 8'b00000000 ;
			15'h00005B9C : data <= 8'b00000000 ;
			15'h00005B9D : data <= 8'b00000000 ;
			15'h00005B9E : data <= 8'b00000000 ;
			15'h00005B9F : data <= 8'b00000000 ;
			15'h00005BA0 : data <= 8'b00000000 ;
			15'h00005BA1 : data <= 8'b00000000 ;
			15'h00005BA2 : data <= 8'b00000000 ;
			15'h00005BA3 : data <= 8'b00000000 ;
			15'h00005BA4 : data <= 8'b00000000 ;
			15'h00005BA5 : data <= 8'b00000000 ;
			15'h00005BA6 : data <= 8'b00000000 ;
			15'h00005BA7 : data <= 8'b00000000 ;
			15'h00005BA8 : data <= 8'b00000000 ;
			15'h00005BA9 : data <= 8'b00000000 ;
			15'h00005BAA : data <= 8'b00000000 ;
			15'h00005BAB : data <= 8'b00000000 ;
			15'h00005BAC : data <= 8'b00000000 ;
			15'h00005BAD : data <= 8'b00000000 ;
			15'h00005BAE : data <= 8'b00000000 ;
			15'h00005BAF : data <= 8'b00000000 ;
			15'h00005BB0 : data <= 8'b00000000 ;
			15'h00005BB1 : data <= 8'b00000000 ;
			15'h00005BB2 : data <= 8'b00000000 ;
			15'h00005BB3 : data <= 8'b00000000 ;
			15'h00005BB4 : data <= 8'b00000000 ;
			15'h00005BB5 : data <= 8'b00000000 ;
			15'h00005BB6 : data <= 8'b00000000 ;
			15'h00005BB7 : data <= 8'b00000000 ;
			15'h00005BB8 : data <= 8'b00000000 ;
			15'h00005BB9 : data <= 8'b00000000 ;
			15'h00005BBA : data <= 8'b00000000 ;
			15'h00005BBB : data <= 8'b00000000 ;
			15'h00005BBC : data <= 8'b00000000 ;
			15'h00005BBD : data <= 8'b00000000 ;
			15'h00005BBE : data <= 8'b00000000 ;
			15'h00005BBF : data <= 8'b00000000 ;
			15'h00005BC0 : data <= 8'b00000000 ;
			15'h00005BC1 : data <= 8'b00000000 ;
			15'h00005BC2 : data <= 8'b00000000 ;
			15'h00005BC3 : data <= 8'b00000000 ;
			15'h00005BC4 : data <= 8'b00000000 ;
			15'h00005BC5 : data <= 8'b00000000 ;
			15'h00005BC6 : data <= 8'b00000000 ;
			15'h00005BC7 : data <= 8'b00000000 ;
			15'h00005BC8 : data <= 8'b00000000 ;
			15'h00005BC9 : data <= 8'b00000000 ;
			15'h00005BCA : data <= 8'b00000000 ;
			15'h00005BCB : data <= 8'b00000000 ;
			15'h00005BCC : data <= 8'b00000000 ;
			15'h00005BCD : data <= 8'b00000000 ;
			15'h00005BCE : data <= 8'b00000000 ;
			15'h00005BCF : data <= 8'b00000000 ;
			15'h00005BD0 : data <= 8'b00000000 ;
			15'h00005BD1 : data <= 8'b00000000 ;
			15'h00005BD2 : data <= 8'b00000000 ;
			15'h00005BD3 : data <= 8'b00000000 ;
			15'h00005BD4 : data <= 8'b00000000 ;
			15'h00005BD5 : data <= 8'b00000000 ;
			15'h00005BD6 : data <= 8'b00000000 ;
			15'h00005BD7 : data <= 8'b00000000 ;
			15'h00005BD8 : data <= 8'b00000000 ;
			15'h00005BD9 : data <= 8'b00000000 ;
			15'h00005BDA : data <= 8'b00000000 ;
			15'h00005BDB : data <= 8'b00000000 ;
			15'h00005BDC : data <= 8'b00000000 ;
			15'h00005BDD : data <= 8'b00000000 ;
			15'h00005BDE : data <= 8'b00000000 ;
			15'h00005BDF : data <= 8'b00000000 ;
			15'h00005BE0 : data <= 8'b00000000 ;
			15'h00005BE1 : data <= 8'b00000000 ;
			15'h00005BE2 : data <= 8'b00000000 ;
			15'h00005BE3 : data <= 8'b00000000 ;
			15'h00005BE4 : data <= 8'b00000000 ;
			15'h00005BE5 : data <= 8'b00000000 ;
			15'h00005BE6 : data <= 8'b00000000 ;
			15'h00005BE7 : data <= 8'b00000000 ;
			15'h00005BE8 : data <= 8'b00000000 ;
			15'h00005BE9 : data <= 8'b00000000 ;
			15'h00005BEA : data <= 8'b00000000 ;
			15'h00005BEB : data <= 8'b00000000 ;
			15'h00005BEC : data <= 8'b00000000 ;
			15'h00005BED : data <= 8'b00000000 ;
			15'h00005BEE : data <= 8'b00000000 ;
			15'h00005BEF : data <= 8'b00000000 ;
			15'h00005BF0 : data <= 8'b00000000 ;
			15'h00005BF1 : data <= 8'b00000000 ;
			15'h00005BF2 : data <= 8'b00000000 ;
			15'h00005BF3 : data <= 8'b00000000 ;
			15'h00005BF4 : data <= 8'b00000000 ;
			15'h00005BF5 : data <= 8'b00000000 ;
			15'h00005BF6 : data <= 8'b00000000 ;
			15'h00005BF7 : data <= 8'b00000000 ;
			15'h00005BF8 : data <= 8'b00000000 ;
			15'h00005BF9 : data <= 8'b00000000 ;
			15'h00005BFA : data <= 8'b00000000 ;
			15'h00005BFB : data <= 8'b00000000 ;
			15'h00005BFC : data <= 8'b00000000 ;
			15'h00005BFD : data <= 8'b00000000 ;
			15'h00005BFE : data <= 8'b00000000 ;
			15'h00005BFF : data <= 8'b00000000 ;
			15'h00005C00 : data <= 8'b00000000 ;
			15'h00005C01 : data <= 8'b00000000 ;
			15'h00005C02 : data <= 8'b00000000 ;
			15'h00005C03 : data <= 8'b00000000 ;
			15'h00005C04 : data <= 8'b00000000 ;
			15'h00005C05 : data <= 8'b00000000 ;
			15'h00005C06 : data <= 8'b00000000 ;
			15'h00005C07 : data <= 8'b00000000 ;
			15'h00005C08 : data <= 8'b00000000 ;
			15'h00005C09 : data <= 8'b00000000 ;
			15'h00005C0A : data <= 8'b00000000 ;
			15'h00005C0B : data <= 8'b00000000 ;
			15'h00005C0C : data <= 8'b00000000 ;
			15'h00005C0D : data <= 8'b00000000 ;
			15'h00005C0E : data <= 8'b00000000 ;
			15'h00005C0F : data <= 8'b00000000 ;
			15'h00005C10 : data <= 8'b00000000 ;
			15'h00005C11 : data <= 8'b00000000 ;
			15'h00005C12 : data <= 8'b00000000 ;
			15'h00005C13 : data <= 8'b00000000 ;
			15'h00005C14 : data <= 8'b00000000 ;
			15'h00005C15 : data <= 8'b00000000 ;
			15'h00005C16 : data <= 8'b00000000 ;
			15'h00005C17 : data <= 8'b00000000 ;
			15'h00005C18 : data <= 8'b00000000 ;
			15'h00005C19 : data <= 8'b00000000 ;
			15'h00005C1A : data <= 8'b00000000 ;
			15'h00005C1B : data <= 8'b00000000 ;
			15'h00005C1C : data <= 8'b00000000 ;
			15'h00005C1D : data <= 8'b00000000 ;
			15'h00005C1E : data <= 8'b00000000 ;
			15'h00005C1F : data <= 8'b00000000 ;
			15'h00005C20 : data <= 8'b00000000 ;
			15'h00005C21 : data <= 8'b00000000 ;
			15'h00005C22 : data <= 8'b00000000 ;
			15'h00005C23 : data <= 8'b00000000 ;
			15'h00005C24 : data <= 8'b00000000 ;
			15'h00005C25 : data <= 8'b00000000 ;
			15'h00005C26 : data <= 8'b00000000 ;
			15'h00005C27 : data <= 8'b00000000 ;
			15'h00005C28 : data <= 8'b00000000 ;
			15'h00005C29 : data <= 8'b00000000 ;
			15'h00005C2A : data <= 8'b00000000 ;
			15'h00005C2B : data <= 8'b00000000 ;
			15'h00005C2C : data <= 8'b00000000 ;
			15'h00005C2D : data <= 8'b00000000 ;
			15'h00005C2E : data <= 8'b00000000 ;
			15'h00005C2F : data <= 8'b00000000 ;
			15'h00005C30 : data <= 8'b00000000 ;
			15'h00005C31 : data <= 8'b00000000 ;
			15'h00005C32 : data <= 8'b00000000 ;
			15'h00005C33 : data <= 8'b00000000 ;
			15'h00005C34 : data <= 8'b00000000 ;
			15'h00005C35 : data <= 8'b00000000 ;
			15'h00005C36 : data <= 8'b00000000 ;
			15'h00005C37 : data <= 8'b00000000 ;
			15'h00005C38 : data <= 8'b00000000 ;
			15'h00005C39 : data <= 8'b00000000 ;
			15'h00005C3A : data <= 8'b00000000 ;
			15'h00005C3B : data <= 8'b00000000 ;
			15'h00005C3C : data <= 8'b00000000 ;
			15'h00005C3D : data <= 8'b00000000 ;
			15'h00005C3E : data <= 8'b00000000 ;
			15'h00005C3F : data <= 8'b00000000 ;
			15'h00005C40 : data <= 8'b00000000 ;
			15'h00005C41 : data <= 8'b00000000 ;
			15'h00005C42 : data <= 8'b00000000 ;
			15'h00005C43 : data <= 8'b00000000 ;
			15'h00005C44 : data <= 8'b00000000 ;
			15'h00005C45 : data <= 8'b00000000 ;
			15'h00005C46 : data <= 8'b00000000 ;
			15'h00005C47 : data <= 8'b00000000 ;
			15'h00005C48 : data <= 8'b00000000 ;
			15'h00005C49 : data <= 8'b00000000 ;
			15'h00005C4A : data <= 8'b00000000 ;
			15'h00005C4B : data <= 8'b00000000 ;
			15'h00005C4C : data <= 8'b00000000 ;
			15'h00005C4D : data <= 8'b00000000 ;
			15'h00005C4E : data <= 8'b00000000 ;
			15'h00005C4F : data <= 8'b00000000 ;
			15'h00005C50 : data <= 8'b00000000 ;
			15'h00005C51 : data <= 8'b00000000 ;
			15'h00005C52 : data <= 8'b00000000 ;
			15'h00005C53 : data <= 8'b00000000 ;
			15'h00005C54 : data <= 8'b00000000 ;
			15'h00005C55 : data <= 8'b00000000 ;
			15'h00005C56 : data <= 8'b00000000 ;
			15'h00005C57 : data <= 8'b00000000 ;
			15'h00005C58 : data <= 8'b00000000 ;
			15'h00005C59 : data <= 8'b00000000 ;
			15'h00005C5A : data <= 8'b00000000 ;
			15'h00005C5B : data <= 8'b00000000 ;
			15'h00005C5C : data <= 8'b00000000 ;
			15'h00005C5D : data <= 8'b00000000 ;
			15'h00005C5E : data <= 8'b00000000 ;
			15'h00005C5F : data <= 8'b00000000 ;
			15'h00005C60 : data <= 8'b00000000 ;
			15'h00005C61 : data <= 8'b00000000 ;
			15'h00005C62 : data <= 8'b00000000 ;
			15'h00005C63 : data <= 8'b00000000 ;
			15'h00005C64 : data <= 8'b00000000 ;
			15'h00005C65 : data <= 8'b00000000 ;
			15'h00005C66 : data <= 8'b00000000 ;
			15'h00005C67 : data <= 8'b00000000 ;
			15'h00005C68 : data <= 8'b00000000 ;
			15'h00005C69 : data <= 8'b00000000 ;
			15'h00005C6A : data <= 8'b00000000 ;
			15'h00005C6B : data <= 8'b00000000 ;
			15'h00005C6C : data <= 8'b00000000 ;
			15'h00005C6D : data <= 8'b00000000 ;
			15'h00005C6E : data <= 8'b00000000 ;
			15'h00005C6F : data <= 8'b00000000 ;
			15'h00005C70 : data <= 8'b00000000 ;
			15'h00005C71 : data <= 8'b00000000 ;
			15'h00005C72 : data <= 8'b00000000 ;
			15'h00005C73 : data <= 8'b00000000 ;
			15'h00005C74 : data <= 8'b00000000 ;
			15'h00005C75 : data <= 8'b00000000 ;
			15'h00005C76 : data <= 8'b00000000 ;
			15'h00005C77 : data <= 8'b00000000 ;
			15'h00005C78 : data <= 8'b00000000 ;
			15'h00005C79 : data <= 8'b00000000 ;
			15'h00005C7A : data <= 8'b00000000 ;
			15'h00005C7B : data <= 8'b00000000 ;
			15'h00005C7C : data <= 8'b00000000 ;
			15'h00005C7D : data <= 8'b00000000 ;
			15'h00005C7E : data <= 8'b00000000 ;
			15'h00005C7F : data <= 8'b00000000 ;
			15'h00005C80 : data <= 8'b00000000 ;
			15'h00005C81 : data <= 8'b00000000 ;
			15'h00005C82 : data <= 8'b00000000 ;
			15'h00005C83 : data <= 8'b00000000 ;
			15'h00005C84 : data <= 8'b00000000 ;
			15'h00005C85 : data <= 8'b00000000 ;
			15'h00005C86 : data <= 8'b00000000 ;
			15'h00005C87 : data <= 8'b00000000 ;
			15'h00005C88 : data <= 8'b00000000 ;
			15'h00005C89 : data <= 8'b00000000 ;
			15'h00005C8A : data <= 8'b00000000 ;
			15'h00005C8B : data <= 8'b00000000 ;
			15'h00005C8C : data <= 8'b00000000 ;
			15'h00005C8D : data <= 8'b00000000 ;
			15'h00005C8E : data <= 8'b00000000 ;
			15'h00005C8F : data <= 8'b00000000 ;
			15'h00005C90 : data <= 8'b00000000 ;
			15'h00005C91 : data <= 8'b00000000 ;
			15'h00005C92 : data <= 8'b00000000 ;
			15'h00005C93 : data <= 8'b00000000 ;
			15'h00005C94 : data <= 8'b00000000 ;
			15'h00005C95 : data <= 8'b00000000 ;
			15'h00005C96 : data <= 8'b00000000 ;
			15'h00005C97 : data <= 8'b00000000 ;
			15'h00005C98 : data <= 8'b00000000 ;
			15'h00005C99 : data <= 8'b00000000 ;
			15'h00005C9A : data <= 8'b00000000 ;
			15'h00005C9B : data <= 8'b00000000 ;
			15'h00005C9C : data <= 8'b00000000 ;
			15'h00005C9D : data <= 8'b00000000 ;
			15'h00005C9E : data <= 8'b00000000 ;
			15'h00005C9F : data <= 8'b00000000 ;
			15'h00005CA0 : data <= 8'b00000000 ;
			15'h00005CA1 : data <= 8'b00000000 ;
			15'h00005CA2 : data <= 8'b00000000 ;
			15'h00005CA3 : data <= 8'b00000000 ;
			15'h00005CA4 : data <= 8'b00000000 ;
			15'h00005CA5 : data <= 8'b00000000 ;
			15'h00005CA6 : data <= 8'b00000000 ;
			15'h00005CA7 : data <= 8'b00000000 ;
			15'h00005CA8 : data <= 8'b00000000 ;
			15'h00005CA9 : data <= 8'b00000000 ;
			15'h00005CAA : data <= 8'b00000000 ;
			15'h00005CAB : data <= 8'b00000000 ;
			15'h00005CAC : data <= 8'b00000000 ;
			15'h00005CAD : data <= 8'b00000000 ;
			15'h00005CAE : data <= 8'b00000000 ;
			15'h00005CAF : data <= 8'b00000000 ;
			15'h00005CB0 : data <= 8'b00000000 ;
			15'h00005CB1 : data <= 8'b00000000 ;
			15'h00005CB2 : data <= 8'b00000000 ;
			15'h00005CB3 : data <= 8'b00000000 ;
			15'h00005CB4 : data <= 8'b00000000 ;
			15'h00005CB5 : data <= 8'b00000000 ;
			15'h00005CB6 : data <= 8'b00000000 ;
			15'h00005CB7 : data <= 8'b00000000 ;
			15'h00005CB8 : data <= 8'b00000000 ;
			15'h00005CB9 : data <= 8'b00000000 ;
			15'h00005CBA : data <= 8'b00000000 ;
			15'h00005CBB : data <= 8'b00000000 ;
			15'h00005CBC : data <= 8'b00000000 ;
			15'h00005CBD : data <= 8'b00000000 ;
			15'h00005CBE : data <= 8'b00000000 ;
			15'h00005CBF : data <= 8'b00000000 ;
			15'h00005CC0 : data <= 8'b00000000 ;
			15'h00005CC1 : data <= 8'b00000000 ;
			15'h00005CC2 : data <= 8'b00000000 ;
			15'h00005CC3 : data <= 8'b00000000 ;
			15'h00005CC4 : data <= 8'b00000000 ;
			15'h00005CC5 : data <= 8'b00000000 ;
			15'h00005CC6 : data <= 8'b00000000 ;
			15'h00005CC7 : data <= 8'b00000000 ;
			15'h00005CC8 : data <= 8'b00000000 ;
			15'h00005CC9 : data <= 8'b00000000 ;
			15'h00005CCA : data <= 8'b00000000 ;
			15'h00005CCB : data <= 8'b00000000 ;
			15'h00005CCC : data <= 8'b00000000 ;
			15'h00005CCD : data <= 8'b00000000 ;
			15'h00005CCE : data <= 8'b00000000 ;
			15'h00005CCF : data <= 8'b00000000 ;
			15'h00005CD0 : data <= 8'b00000000 ;
			15'h00005CD1 : data <= 8'b00000000 ;
			15'h00005CD2 : data <= 8'b00000000 ;
			15'h00005CD3 : data <= 8'b00000000 ;
			15'h00005CD4 : data <= 8'b00000000 ;
			15'h00005CD5 : data <= 8'b00000000 ;
			15'h00005CD6 : data <= 8'b00000000 ;
			15'h00005CD7 : data <= 8'b00000000 ;
			15'h00005CD8 : data <= 8'b00000000 ;
			15'h00005CD9 : data <= 8'b00000000 ;
			15'h00005CDA : data <= 8'b00000000 ;
			15'h00005CDB : data <= 8'b00000000 ;
			15'h00005CDC : data <= 8'b00000000 ;
			15'h00005CDD : data <= 8'b00000000 ;
			15'h00005CDE : data <= 8'b00000000 ;
			15'h00005CDF : data <= 8'b00000000 ;
			15'h00005CE0 : data <= 8'b00000000 ;
			15'h00005CE1 : data <= 8'b00000000 ;
			15'h00005CE2 : data <= 8'b00000000 ;
			15'h00005CE3 : data <= 8'b00000000 ;
			15'h00005CE4 : data <= 8'b00000000 ;
			15'h00005CE5 : data <= 8'b00000000 ;
			15'h00005CE6 : data <= 8'b00000000 ;
			15'h00005CE7 : data <= 8'b00000000 ;
			15'h00005CE8 : data <= 8'b00000000 ;
			15'h00005CE9 : data <= 8'b00000000 ;
			15'h00005CEA : data <= 8'b00000000 ;
			15'h00005CEB : data <= 8'b00000000 ;
			15'h00005CEC : data <= 8'b00000000 ;
			15'h00005CED : data <= 8'b00000000 ;
			15'h00005CEE : data <= 8'b00000000 ;
			15'h00005CEF : data <= 8'b00000000 ;
			15'h00005CF0 : data <= 8'b00000000 ;
			15'h00005CF1 : data <= 8'b00000000 ;
			15'h00005CF2 : data <= 8'b00000000 ;
			15'h00005CF3 : data <= 8'b00000000 ;
			15'h00005CF4 : data <= 8'b00000000 ;
			15'h00005CF5 : data <= 8'b00000000 ;
			15'h00005CF6 : data <= 8'b00000000 ;
			15'h00005CF7 : data <= 8'b00000000 ;
			15'h00005CF8 : data <= 8'b00000000 ;
			15'h00005CF9 : data <= 8'b00000000 ;
			15'h00005CFA : data <= 8'b00000000 ;
			15'h00005CFB : data <= 8'b00000000 ;
			15'h00005CFC : data <= 8'b00000000 ;
			15'h00005CFD : data <= 8'b00000000 ;
			15'h00005CFE : data <= 8'b00000000 ;
			15'h00005CFF : data <= 8'b00000000 ;
			15'h00005D00 : data <= 8'b00000000 ;
			15'h00005D01 : data <= 8'b00000000 ;
			15'h00005D02 : data <= 8'b00000000 ;
			15'h00005D03 : data <= 8'b00000000 ;
			15'h00005D04 : data <= 8'b00000000 ;
			15'h00005D05 : data <= 8'b00000000 ;
			15'h00005D06 : data <= 8'b00000000 ;
			15'h00005D07 : data <= 8'b00000000 ;
			15'h00005D08 : data <= 8'b00000000 ;
			15'h00005D09 : data <= 8'b00000000 ;
			15'h00005D0A : data <= 8'b00000000 ;
			15'h00005D0B : data <= 8'b00000000 ;
			15'h00005D0C : data <= 8'b00000000 ;
			15'h00005D0D : data <= 8'b00000000 ;
			15'h00005D0E : data <= 8'b00000000 ;
			15'h00005D0F : data <= 8'b00000000 ;
			15'h00005D10 : data <= 8'b00000000 ;
			15'h00005D11 : data <= 8'b00000000 ;
			15'h00005D12 : data <= 8'b00000000 ;
			15'h00005D13 : data <= 8'b00000000 ;
			15'h00005D14 : data <= 8'b00000000 ;
			15'h00005D15 : data <= 8'b00000000 ;
			15'h00005D16 : data <= 8'b00000000 ;
			15'h00005D17 : data <= 8'b00000000 ;
			15'h00005D18 : data <= 8'b00000000 ;
			15'h00005D19 : data <= 8'b00000000 ;
			15'h00005D1A : data <= 8'b00000000 ;
			15'h00005D1B : data <= 8'b00000000 ;
			15'h00005D1C : data <= 8'b00000000 ;
			15'h00005D1D : data <= 8'b00000000 ;
			15'h00005D1E : data <= 8'b00000000 ;
			15'h00005D1F : data <= 8'b00000000 ;
			15'h00005D20 : data <= 8'b00000000 ;
			15'h00005D21 : data <= 8'b00000000 ;
			15'h00005D22 : data <= 8'b00000000 ;
			15'h00005D23 : data <= 8'b00000000 ;
			15'h00005D24 : data <= 8'b00000000 ;
			15'h00005D25 : data <= 8'b00000000 ;
			15'h00005D26 : data <= 8'b00000000 ;
			15'h00005D27 : data <= 8'b00000000 ;
			15'h00005D28 : data <= 8'b00000000 ;
			15'h00005D29 : data <= 8'b00000000 ;
			15'h00005D2A : data <= 8'b00000000 ;
			15'h00005D2B : data <= 8'b00000000 ;
			15'h00005D2C : data <= 8'b00000000 ;
			15'h00005D2D : data <= 8'b00000000 ;
			15'h00005D2E : data <= 8'b00000000 ;
			15'h00005D2F : data <= 8'b00000000 ;
			15'h00005D30 : data <= 8'b00000000 ;
			15'h00005D31 : data <= 8'b00000000 ;
			15'h00005D32 : data <= 8'b00000000 ;
			15'h00005D33 : data <= 8'b00000000 ;
			15'h00005D34 : data <= 8'b00000000 ;
			15'h00005D35 : data <= 8'b00000000 ;
			15'h00005D36 : data <= 8'b00000000 ;
			15'h00005D37 : data <= 8'b00000000 ;
			15'h00005D38 : data <= 8'b00000000 ;
			15'h00005D39 : data <= 8'b00000000 ;
			15'h00005D3A : data <= 8'b00000000 ;
			15'h00005D3B : data <= 8'b00000000 ;
			15'h00005D3C : data <= 8'b00000000 ;
			15'h00005D3D : data <= 8'b00000000 ;
			15'h00005D3E : data <= 8'b00000000 ;
			15'h00005D3F : data <= 8'b00000000 ;
			15'h00005D40 : data <= 8'b00000000 ;
			15'h00005D41 : data <= 8'b00000000 ;
			15'h00005D42 : data <= 8'b00000000 ;
			15'h00005D43 : data <= 8'b00000000 ;
			15'h00005D44 : data <= 8'b00000000 ;
			15'h00005D45 : data <= 8'b00000000 ;
			15'h00005D46 : data <= 8'b00000000 ;
			15'h00005D47 : data <= 8'b00000000 ;
			15'h00005D48 : data <= 8'b00000000 ;
			15'h00005D49 : data <= 8'b00000000 ;
			15'h00005D4A : data <= 8'b00000000 ;
			15'h00005D4B : data <= 8'b00000000 ;
			15'h00005D4C : data <= 8'b00000000 ;
			15'h00005D4D : data <= 8'b00000000 ;
			15'h00005D4E : data <= 8'b00000000 ;
			15'h00005D4F : data <= 8'b00000000 ;
			15'h00005D50 : data <= 8'b00000000 ;
			15'h00005D51 : data <= 8'b00000000 ;
			15'h00005D52 : data <= 8'b00000000 ;
			15'h00005D53 : data <= 8'b00000000 ;
			15'h00005D54 : data <= 8'b00000000 ;
			15'h00005D55 : data <= 8'b00000000 ;
			15'h00005D56 : data <= 8'b00000000 ;
			15'h00005D57 : data <= 8'b00000000 ;
			15'h00005D58 : data <= 8'b00000000 ;
			15'h00005D59 : data <= 8'b00000000 ;
			15'h00005D5A : data <= 8'b00000000 ;
			15'h00005D5B : data <= 8'b00000000 ;
			15'h00005D5C : data <= 8'b00000000 ;
			15'h00005D5D : data <= 8'b00000000 ;
			15'h00005D5E : data <= 8'b00000000 ;
			15'h00005D5F : data <= 8'b00000000 ;
			15'h00005D60 : data <= 8'b00000000 ;
			15'h00005D61 : data <= 8'b00000000 ;
			15'h00005D62 : data <= 8'b00000000 ;
			15'h00005D63 : data <= 8'b00000000 ;
			15'h00005D64 : data <= 8'b00000000 ;
			15'h00005D65 : data <= 8'b00000000 ;
			15'h00005D66 : data <= 8'b00000000 ;
			15'h00005D67 : data <= 8'b00000000 ;
			15'h00005D68 : data <= 8'b00000000 ;
			15'h00005D69 : data <= 8'b00000000 ;
			15'h00005D6A : data <= 8'b00000000 ;
			15'h00005D6B : data <= 8'b00000000 ;
			15'h00005D6C : data <= 8'b00000000 ;
			15'h00005D6D : data <= 8'b00000000 ;
			15'h00005D6E : data <= 8'b00000000 ;
			15'h00005D6F : data <= 8'b00000000 ;
			15'h00005D70 : data <= 8'b00000000 ;
			15'h00005D71 : data <= 8'b00000000 ;
			15'h00005D72 : data <= 8'b00000000 ;
			15'h00005D73 : data <= 8'b00000000 ;
			15'h00005D74 : data <= 8'b00000000 ;
			15'h00005D75 : data <= 8'b00000000 ;
			15'h00005D76 : data <= 8'b00000000 ;
			15'h00005D77 : data <= 8'b00000000 ;
			15'h00005D78 : data <= 8'b00000000 ;
			15'h00005D79 : data <= 8'b00000000 ;
			15'h00005D7A : data <= 8'b00000000 ;
			15'h00005D7B : data <= 8'b00000000 ;
			15'h00005D7C : data <= 8'b00000000 ;
			15'h00005D7D : data <= 8'b00000000 ;
			15'h00005D7E : data <= 8'b00000000 ;
			15'h00005D7F : data <= 8'b00000000 ;
			15'h00005D80 : data <= 8'b00000000 ;
			15'h00005D81 : data <= 8'b00000000 ;
			15'h00005D82 : data <= 8'b00000000 ;
			15'h00005D83 : data <= 8'b00000000 ;
			15'h00005D84 : data <= 8'b00000000 ;
			15'h00005D85 : data <= 8'b00000000 ;
			15'h00005D86 : data <= 8'b00000000 ;
			15'h00005D87 : data <= 8'b00000000 ;
			15'h00005D88 : data <= 8'b00000000 ;
			15'h00005D89 : data <= 8'b00000000 ;
			15'h00005D8A : data <= 8'b00000000 ;
			15'h00005D8B : data <= 8'b00000000 ;
			15'h00005D8C : data <= 8'b00000000 ;
			15'h00005D8D : data <= 8'b00000000 ;
			15'h00005D8E : data <= 8'b00000000 ;
			15'h00005D8F : data <= 8'b00000000 ;
			15'h00005D90 : data <= 8'b00000000 ;
			15'h00005D91 : data <= 8'b00000000 ;
			15'h00005D92 : data <= 8'b00000000 ;
			15'h00005D93 : data <= 8'b00000000 ;
			15'h00005D94 : data <= 8'b00000000 ;
			15'h00005D95 : data <= 8'b00000000 ;
			15'h00005D96 : data <= 8'b00000000 ;
			15'h00005D97 : data <= 8'b00000000 ;
			15'h00005D98 : data <= 8'b00000000 ;
			15'h00005D99 : data <= 8'b00000000 ;
			15'h00005D9A : data <= 8'b00000000 ;
			15'h00005D9B : data <= 8'b00000000 ;
			15'h00005D9C : data <= 8'b00000000 ;
			15'h00005D9D : data <= 8'b00000000 ;
			15'h00005D9E : data <= 8'b00000000 ;
			15'h00005D9F : data <= 8'b00000000 ;
			15'h00005DA0 : data <= 8'b00000000 ;
			15'h00005DA1 : data <= 8'b00000000 ;
			15'h00005DA2 : data <= 8'b00000000 ;
			15'h00005DA3 : data <= 8'b00000000 ;
			15'h00005DA4 : data <= 8'b00000000 ;
			15'h00005DA5 : data <= 8'b00000000 ;
			15'h00005DA6 : data <= 8'b00000000 ;
			15'h00005DA7 : data <= 8'b00000000 ;
			15'h00005DA8 : data <= 8'b00000000 ;
			15'h00005DA9 : data <= 8'b00000000 ;
			15'h00005DAA : data <= 8'b00000000 ;
			15'h00005DAB : data <= 8'b00000000 ;
			15'h00005DAC : data <= 8'b00000000 ;
			15'h00005DAD : data <= 8'b00000000 ;
			15'h00005DAE : data <= 8'b00000000 ;
			15'h00005DAF : data <= 8'b00000000 ;
			15'h00005DB0 : data <= 8'b00000000 ;
			15'h00005DB1 : data <= 8'b00000000 ;
			15'h00005DB2 : data <= 8'b00000000 ;
			15'h00005DB3 : data <= 8'b00000000 ;
			15'h00005DB4 : data <= 8'b00000000 ;
			15'h00005DB5 : data <= 8'b00000000 ;
			15'h00005DB6 : data <= 8'b00000000 ;
			15'h00005DB7 : data <= 8'b00000000 ;
			15'h00005DB8 : data <= 8'b00000000 ;
			15'h00005DB9 : data <= 8'b00000000 ;
			15'h00005DBA : data <= 8'b00000000 ;
			15'h00005DBB : data <= 8'b00000000 ;
			15'h00005DBC : data <= 8'b00000000 ;
			15'h00005DBD : data <= 8'b00000000 ;
			15'h00005DBE : data <= 8'b00000000 ;
			15'h00005DBF : data <= 8'b00000000 ;
			15'h00005DC0 : data <= 8'b00000000 ;
			15'h00005DC1 : data <= 8'b00000000 ;
			15'h00005DC2 : data <= 8'b00000000 ;
			15'h00005DC3 : data <= 8'b00000000 ;
			15'h00005DC4 : data <= 8'b00000000 ;
			15'h00005DC5 : data <= 8'b00000000 ;
			15'h00005DC6 : data <= 8'b00000000 ;
			15'h00005DC7 : data <= 8'b00000000 ;
			15'h00005DC8 : data <= 8'b00000000 ;
			15'h00005DC9 : data <= 8'b00000000 ;
			15'h00005DCA : data <= 8'b00000000 ;
			15'h00005DCB : data <= 8'b00000000 ;
			15'h00005DCC : data <= 8'b00000000 ;
			15'h00005DCD : data <= 8'b00000000 ;
			15'h00005DCE : data <= 8'b00000000 ;
			15'h00005DCF : data <= 8'b00000000 ;
			15'h00005DD0 : data <= 8'b00000000 ;
			15'h00005DD1 : data <= 8'b00000000 ;
			15'h00005DD2 : data <= 8'b00000000 ;
			15'h00005DD3 : data <= 8'b00000000 ;
			15'h00005DD4 : data <= 8'b00000000 ;
			15'h00005DD5 : data <= 8'b00000000 ;
			15'h00005DD6 : data <= 8'b00000000 ;
			15'h00005DD7 : data <= 8'b00000000 ;
			15'h00005DD8 : data <= 8'b00000000 ;
			15'h00005DD9 : data <= 8'b00000000 ;
			15'h00005DDA : data <= 8'b00000000 ;
			15'h00005DDB : data <= 8'b00000000 ;
			15'h00005DDC : data <= 8'b00000000 ;
			15'h00005DDD : data <= 8'b00000000 ;
			15'h00005DDE : data <= 8'b00000000 ;
			15'h00005DDF : data <= 8'b00000000 ;
			15'h00005DE0 : data <= 8'b00000000 ;
			15'h00005DE1 : data <= 8'b00000000 ;
			15'h00005DE2 : data <= 8'b00000000 ;
			15'h00005DE3 : data <= 8'b00000000 ;
			15'h00005DE4 : data <= 8'b00000000 ;
			15'h00005DE5 : data <= 8'b00000000 ;
			15'h00005DE6 : data <= 8'b00000000 ;
			15'h00005DE7 : data <= 8'b00000000 ;
			15'h00005DE8 : data <= 8'b00000000 ;
			15'h00005DE9 : data <= 8'b00000000 ;
			15'h00005DEA : data <= 8'b00000000 ;
			15'h00005DEB : data <= 8'b00000000 ;
			15'h00005DEC : data <= 8'b00000000 ;
			15'h00005DED : data <= 8'b00000000 ;
			15'h00005DEE : data <= 8'b00000000 ;
			15'h00005DEF : data <= 8'b00000000 ;
			15'h00005DF0 : data <= 8'b00000000 ;
			15'h00005DF1 : data <= 8'b00000000 ;
			15'h00005DF2 : data <= 8'b00000000 ;
			15'h00005DF3 : data <= 8'b00000000 ;
			15'h00005DF4 : data <= 8'b00000000 ;
			15'h00005DF5 : data <= 8'b00000000 ;
			15'h00005DF6 : data <= 8'b00000000 ;
			15'h00005DF7 : data <= 8'b00000000 ;
			15'h00005DF8 : data <= 8'b00000000 ;
			15'h00005DF9 : data <= 8'b00000000 ;
			15'h00005DFA : data <= 8'b00000000 ;
			15'h00005DFB : data <= 8'b00000000 ;
			15'h00005DFC : data <= 8'b00000000 ;
			15'h00005DFD : data <= 8'b00000000 ;
			15'h00005DFE : data <= 8'b00000000 ;
			15'h00005DFF : data <= 8'b00000000 ;
			15'h00005E00 : data <= 8'b00000000 ;
			15'h00005E01 : data <= 8'b00000000 ;
			15'h00005E02 : data <= 8'b00000000 ;
			15'h00005E03 : data <= 8'b00000000 ;
			15'h00005E04 : data <= 8'b00000000 ;
			15'h00005E05 : data <= 8'b00000000 ;
			15'h00005E06 : data <= 8'b00000000 ;
			15'h00005E07 : data <= 8'b00000000 ;
			15'h00005E08 : data <= 8'b00000000 ;
			15'h00005E09 : data <= 8'b00000000 ;
			15'h00005E0A : data <= 8'b00000000 ;
			15'h00005E0B : data <= 8'b00000000 ;
			15'h00005E0C : data <= 8'b00000000 ;
			15'h00005E0D : data <= 8'b00000000 ;
			15'h00005E0E : data <= 8'b00000000 ;
			15'h00005E0F : data <= 8'b00000000 ;
			15'h00005E10 : data <= 8'b00000000 ;
			15'h00005E11 : data <= 8'b00000000 ;
			15'h00005E12 : data <= 8'b00000000 ;
			15'h00005E13 : data <= 8'b00000000 ;
			15'h00005E14 : data <= 8'b00000000 ;
			15'h00005E15 : data <= 8'b00000000 ;
			15'h00005E16 : data <= 8'b00000000 ;
			15'h00005E17 : data <= 8'b00000000 ;
			15'h00005E18 : data <= 8'b00000000 ;
			15'h00005E19 : data <= 8'b00000000 ;
			15'h00005E1A : data <= 8'b00000000 ;
			15'h00005E1B : data <= 8'b00000000 ;
			15'h00005E1C : data <= 8'b00000000 ;
			15'h00005E1D : data <= 8'b00000000 ;
			15'h00005E1E : data <= 8'b00000000 ;
			15'h00005E1F : data <= 8'b00000000 ;
			15'h00005E20 : data <= 8'b00000000 ;
			15'h00005E21 : data <= 8'b00000000 ;
			15'h00005E22 : data <= 8'b00000000 ;
			15'h00005E23 : data <= 8'b00000000 ;
			15'h00005E24 : data <= 8'b00000000 ;
			15'h00005E25 : data <= 8'b00000000 ;
			15'h00005E26 : data <= 8'b00000000 ;
			15'h00005E27 : data <= 8'b00000000 ;
			15'h00005E28 : data <= 8'b00000000 ;
			15'h00005E29 : data <= 8'b00000000 ;
			15'h00005E2A : data <= 8'b00000000 ;
			15'h00005E2B : data <= 8'b00000000 ;
			15'h00005E2C : data <= 8'b00000000 ;
			15'h00005E2D : data <= 8'b00000000 ;
			15'h00005E2E : data <= 8'b00000000 ;
			15'h00005E2F : data <= 8'b00000000 ;
			15'h00005E30 : data <= 8'b00000000 ;
			15'h00005E31 : data <= 8'b00000000 ;
			15'h00005E32 : data <= 8'b00000000 ;
			15'h00005E33 : data <= 8'b00000000 ;
			15'h00005E34 : data <= 8'b00000000 ;
			15'h00005E35 : data <= 8'b00000000 ;
			15'h00005E36 : data <= 8'b00000000 ;
			15'h00005E37 : data <= 8'b00000000 ;
			15'h00005E38 : data <= 8'b00000000 ;
			15'h00005E39 : data <= 8'b00000000 ;
			15'h00005E3A : data <= 8'b00000000 ;
			15'h00005E3B : data <= 8'b00000000 ;
			15'h00005E3C : data <= 8'b00000000 ;
			15'h00005E3D : data <= 8'b00000000 ;
			15'h00005E3E : data <= 8'b00000000 ;
			15'h00005E3F : data <= 8'b00000000 ;
			15'h00005E40 : data <= 8'b00000000 ;
			15'h00005E41 : data <= 8'b00000000 ;
			15'h00005E42 : data <= 8'b00000000 ;
			15'h00005E43 : data <= 8'b00000000 ;
			15'h00005E44 : data <= 8'b00000000 ;
			15'h00005E45 : data <= 8'b00000000 ;
			15'h00005E46 : data <= 8'b00000000 ;
			15'h00005E47 : data <= 8'b00000000 ;
			15'h00005E48 : data <= 8'b00000000 ;
			15'h00005E49 : data <= 8'b00000000 ;
			15'h00005E4A : data <= 8'b00000000 ;
			15'h00005E4B : data <= 8'b00000000 ;
			15'h00005E4C : data <= 8'b00000000 ;
			15'h00005E4D : data <= 8'b00000000 ;
			15'h00005E4E : data <= 8'b00000000 ;
			15'h00005E4F : data <= 8'b00000000 ;
			15'h00005E50 : data <= 8'b00000000 ;
			15'h00005E51 : data <= 8'b00000000 ;
			15'h00005E52 : data <= 8'b00000000 ;
			15'h00005E53 : data <= 8'b00000000 ;
			15'h00005E54 : data <= 8'b00000000 ;
			15'h00005E55 : data <= 8'b00000000 ;
			15'h00005E56 : data <= 8'b00000000 ;
			15'h00005E57 : data <= 8'b00000000 ;
			15'h00005E58 : data <= 8'b00000000 ;
			15'h00005E59 : data <= 8'b00000000 ;
			15'h00005E5A : data <= 8'b00000000 ;
			15'h00005E5B : data <= 8'b00000000 ;
			15'h00005E5C : data <= 8'b00000000 ;
			15'h00005E5D : data <= 8'b00000000 ;
			15'h00005E5E : data <= 8'b00000000 ;
			15'h00005E5F : data <= 8'b00000000 ;
			15'h00005E60 : data <= 8'b00000000 ;
			15'h00005E61 : data <= 8'b00000000 ;
			15'h00005E62 : data <= 8'b00000000 ;
			15'h00005E63 : data <= 8'b00000000 ;
			15'h00005E64 : data <= 8'b00000000 ;
			15'h00005E65 : data <= 8'b00000000 ;
			15'h00005E66 : data <= 8'b00000000 ;
			15'h00005E67 : data <= 8'b00000000 ;
			15'h00005E68 : data <= 8'b00000000 ;
			15'h00005E69 : data <= 8'b00000000 ;
			15'h00005E6A : data <= 8'b00000000 ;
			15'h00005E6B : data <= 8'b00000000 ;
			15'h00005E6C : data <= 8'b00000000 ;
			15'h00005E6D : data <= 8'b00000000 ;
			15'h00005E6E : data <= 8'b00000000 ;
			15'h00005E6F : data <= 8'b00000000 ;
			15'h00005E70 : data <= 8'b00000000 ;
			15'h00005E71 : data <= 8'b00000000 ;
			15'h00005E72 : data <= 8'b00000000 ;
			15'h00005E73 : data <= 8'b00000000 ;
			15'h00005E74 : data <= 8'b00000000 ;
			15'h00005E75 : data <= 8'b00000000 ;
			15'h00005E76 : data <= 8'b00000000 ;
			15'h00005E77 : data <= 8'b00000000 ;
			15'h00005E78 : data <= 8'b00000000 ;
			15'h00005E79 : data <= 8'b00000000 ;
			15'h00005E7A : data <= 8'b00000000 ;
			15'h00005E7B : data <= 8'b00000000 ;
			15'h00005E7C : data <= 8'b00000000 ;
			15'h00005E7D : data <= 8'b00000000 ;
			15'h00005E7E : data <= 8'b00000000 ;
			15'h00005E7F : data <= 8'b00000000 ;
			15'h00005E80 : data <= 8'b00000000 ;
			15'h00005E81 : data <= 8'b00000000 ;
			15'h00005E82 : data <= 8'b00000000 ;
			15'h00005E83 : data <= 8'b00000000 ;
			15'h00005E84 : data <= 8'b00000000 ;
			15'h00005E85 : data <= 8'b00000000 ;
			15'h00005E86 : data <= 8'b00000000 ;
			15'h00005E87 : data <= 8'b00000000 ;
			15'h00005E88 : data <= 8'b00000000 ;
			15'h00005E89 : data <= 8'b00000000 ;
			15'h00005E8A : data <= 8'b00000000 ;
			15'h00005E8B : data <= 8'b00000000 ;
			15'h00005E8C : data <= 8'b00000000 ;
			15'h00005E8D : data <= 8'b00000000 ;
			15'h00005E8E : data <= 8'b00000000 ;
			15'h00005E8F : data <= 8'b00000000 ;
			15'h00005E90 : data <= 8'b00000000 ;
			15'h00005E91 : data <= 8'b00000000 ;
			15'h00005E92 : data <= 8'b00000000 ;
			15'h00005E93 : data <= 8'b00000000 ;
			15'h00005E94 : data <= 8'b00000000 ;
			15'h00005E95 : data <= 8'b00000000 ;
			15'h00005E96 : data <= 8'b00000000 ;
			15'h00005E97 : data <= 8'b00000000 ;
			15'h00005E98 : data <= 8'b00000000 ;
			15'h00005E99 : data <= 8'b00000000 ;
			15'h00005E9A : data <= 8'b00000000 ;
			15'h00005E9B : data <= 8'b00000000 ;
			15'h00005E9C : data <= 8'b00000000 ;
			15'h00005E9D : data <= 8'b00000000 ;
			15'h00005E9E : data <= 8'b00000000 ;
			15'h00005E9F : data <= 8'b00000000 ;
			15'h00005EA0 : data <= 8'b00000000 ;
			15'h00005EA1 : data <= 8'b00000000 ;
			15'h00005EA2 : data <= 8'b00000000 ;
			15'h00005EA3 : data <= 8'b00000000 ;
			15'h00005EA4 : data <= 8'b00000000 ;
			15'h00005EA5 : data <= 8'b00000000 ;
			15'h00005EA6 : data <= 8'b00000000 ;
			15'h00005EA7 : data <= 8'b00000000 ;
			15'h00005EA8 : data <= 8'b00000000 ;
			15'h00005EA9 : data <= 8'b00000000 ;
			15'h00005EAA : data <= 8'b00000000 ;
			15'h00005EAB : data <= 8'b00000000 ;
			15'h00005EAC : data <= 8'b00000000 ;
			15'h00005EAD : data <= 8'b00000000 ;
			15'h00005EAE : data <= 8'b00000000 ;
			15'h00005EAF : data <= 8'b00000000 ;
			15'h00005EB0 : data <= 8'b00000000 ;
			15'h00005EB1 : data <= 8'b00000000 ;
			15'h00005EB2 : data <= 8'b00000000 ;
			15'h00005EB3 : data <= 8'b00000000 ;
			15'h00005EB4 : data <= 8'b00000000 ;
			15'h00005EB5 : data <= 8'b00000000 ;
			15'h00005EB6 : data <= 8'b00000000 ;
			15'h00005EB7 : data <= 8'b00000000 ;
			15'h00005EB8 : data <= 8'b00000000 ;
			15'h00005EB9 : data <= 8'b00000000 ;
			15'h00005EBA : data <= 8'b00000000 ;
			15'h00005EBB : data <= 8'b00000000 ;
			15'h00005EBC : data <= 8'b00000000 ;
			15'h00005EBD : data <= 8'b00000000 ;
			15'h00005EBE : data <= 8'b00000000 ;
			15'h00005EBF : data <= 8'b00000000 ;
			15'h00005EC0 : data <= 8'b00000000 ;
			15'h00005EC1 : data <= 8'b00000000 ;
			15'h00005EC2 : data <= 8'b00000000 ;
			15'h00005EC3 : data <= 8'b00000000 ;
			15'h00005EC4 : data <= 8'b00000000 ;
			15'h00005EC5 : data <= 8'b00000000 ;
			15'h00005EC6 : data <= 8'b00000000 ;
			15'h00005EC7 : data <= 8'b00000000 ;
			15'h00005EC8 : data <= 8'b00000000 ;
			15'h00005EC9 : data <= 8'b00000000 ;
			15'h00005ECA : data <= 8'b00000000 ;
			15'h00005ECB : data <= 8'b00000000 ;
			15'h00005ECC : data <= 8'b00000000 ;
			15'h00005ECD : data <= 8'b00000000 ;
			15'h00005ECE : data <= 8'b00000000 ;
			15'h00005ECF : data <= 8'b00000000 ;
			15'h00005ED0 : data <= 8'b00000000 ;
			15'h00005ED1 : data <= 8'b00000000 ;
			15'h00005ED2 : data <= 8'b00000000 ;
			15'h00005ED3 : data <= 8'b00000000 ;
			15'h00005ED4 : data <= 8'b00000000 ;
			15'h00005ED5 : data <= 8'b00000000 ;
			15'h00005ED6 : data <= 8'b00000000 ;
			15'h00005ED7 : data <= 8'b00000000 ;
			15'h00005ED8 : data <= 8'b00000000 ;
			15'h00005ED9 : data <= 8'b00000000 ;
			15'h00005EDA : data <= 8'b00000000 ;
			15'h00005EDB : data <= 8'b00000000 ;
			15'h00005EDC : data <= 8'b00000000 ;
			15'h00005EDD : data <= 8'b00000000 ;
			15'h00005EDE : data <= 8'b00000000 ;
			15'h00005EDF : data <= 8'b00000000 ;
			15'h00005EE0 : data <= 8'b00000000 ;
			15'h00005EE1 : data <= 8'b00000000 ;
			15'h00005EE2 : data <= 8'b00000000 ;
			15'h00005EE3 : data <= 8'b00000000 ;
			15'h00005EE4 : data <= 8'b00000000 ;
			15'h00005EE5 : data <= 8'b00000000 ;
			15'h00005EE6 : data <= 8'b00000000 ;
			15'h00005EE7 : data <= 8'b00000000 ;
			15'h00005EE8 : data <= 8'b00000000 ;
			15'h00005EE9 : data <= 8'b00000000 ;
			15'h00005EEA : data <= 8'b00000000 ;
			15'h00005EEB : data <= 8'b00000000 ;
			15'h00005EEC : data <= 8'b00000000 ;
			15'h00005EED : data <= 8'b00000000 ;
			15'h00005EEE : data <= 8'b00000000 ;
			15'h00005EEF : data <= 8'b00000000 ;
			15'h00005EF0 : data <= 8'b00000000 ;
			15'h00005EF1 : data <= 8'b00000000 ;
			15'h00005EF2 : data <= 8'b00000000 ;
			15'h00005EF3 : data <= 8'b00000000 ;
			15'h00005EF4 : data <= 8'b00000000 ;
			15'h00005EF5 : data <= 8'b00000000 ;
			15'h00005EF6 : data <= 8'b00000000 ;
			15'h00005EF7 : data <= 8'b00000000 ;
			15'h00005EF8 : data <= 8'b00000000 ;
			15'h00005EF9 : data <= 8'b00000000 ;
			15'h00005EFA : data <= 8'b00000000 ;
			15'h00005EFB : data <= 8'b00000000 ;
			15'h00005EFC : data <= 8'b00000000 ;
			15'h00005EFD : data <= 8'b00000000 ;
			15'h00005EFE : data <= 8'b00000000 ;
			15'h00005EFF : data <= 8'b00000000 ;
			15'h00005F00 : data <= 8'b00000000 ;
			15'h00005F01 : data <= 8'b00000000 ;
			15'h00005F02 : data <= 8'b00000000 ;
			15'h00005F03 : data <= 8'b00000000 ;
			15'h00005F04 : data <= 8'b00000000 ;
			15'h00005F05 : data <= 8'b00000000 ;
			15'h00005F06 : data <= 8'b00000000 ;
			15'h00005F07 : data <= 8'b00000000 ;
			15'h00005F08 : data <= 8'b00000000 ;
			15'h00005F09 : data <= 8'b00000000 ;
			15'h00005F0A : data <= 8'b00000000 ;
			15'h00005F0B : data <= 8'b00000000 ;
			15'h00005F0C : data <= 8'b00000000 ;
			15'h00005F0D : data <= 8'b00000000 ;
			15'h00005F0E : data <= 8'b00000000 ;
			15'h00005F0F : data <= 8'b00000000 ;
			15'h00005F10 : data <= 8'b00000000 ;
			15'h00005F11 : data <= 8'b00000000 ;
			15'h00005F12 : data <= 8'b00000000 ;
			15'h00005F13 : data <= 8'b00000000 ;
			15'h00005F14 : data <= 8'b00000000 ;
			15'h00005F15 : data <= 8'b00000000 ;
			15'h00005F16 : data <= 8'b00000000 ;
			15'h00005F17 : data <= 8'b00000000 ;
			15'h00005F18 : data <= 8'b00000000 ;
			15'h00005F19 : data <= 8'b00000000 ;
			15'h00005F1A : data <= 8'b00000000 ;
			15'h00005F1B : data <= 8'b00000000 ;
			15'h00005F1C : data <= 8'b00000000 ;
			15'h00005F1D : data <= 8'b00000000 ;
			15'h00005F1E : data <= 8'b00000000 ;
			15'h00005F1F : data <= 8'b00000000 ;
			15'h00005F20 : data <= 8'b00000000 ;
			15'h00005F21 : data <= 8'b00000000 ;
			15'h00005F22 : data <= 8'b00000000 ;
			15'h00005F23 : data <= 8'b00000000 ;
			15'h00005F24 : data <= 8'b00000000 ;
			15'h00005F25 : data <= 8'b00000000 ;
			15'h00005F26 : data <= 8'b00000000 ;
			15'h00005F27 : data <= 8'b00000000 ;
			15'h00005F28 : data <= 8'b00000000 ;
			15'h00005F29 : data <= 8'b00000000 ;
			15'h00005F2A : data <= 8'b00000000 ;
			15'h00005F2B : data <= 8'b00000000 ;
			15'h00005F2C : data <= 8'b00000000 ;
			15'h00005F2D : data <= 8'b00000000 ;
			15'h00005F2E : data <= 8'b00000000 ;
			15'h00005F2F : data <= 8'b00000000 ;
			15'h00005F30 : data <= 8'b00000000 ;
			15'h00005F31 : data <= 8'b00000000 ;
			15'h00005F32 : data <= 8'b00000000 ;
			15'h00005F33 : data <= 8'b00000000 ;
			15'h00005F34 : data <= 8'b00000000 ;
			15'h00005F35 : data <= 8'b00000000 ;
			15'h00005F36 : data <= 8'b00000000 ;
			15'h00005F37 : data <= 8'b00000000 ;
			15'h00005F38 : data <= 8'b00000000 ;
			15'h00005F39 : data <= 8'b00000000 ;
			15'h00005F3A : data <= 8'b00000000 ;
			15'h00005F3B : data <= 8'b00000000 ;
			15'h00005F3C : data <= 8'b00000000 ;
			15'h00005F3D : data <= 8'b00000000 ;
			15'h00005F3E : data <= 8'b00000000 ;
			15'h00005F3F : data <= 8'b00000000 ;
			15'h00005F40 : data <= 8'b00000000 ;
			15'h00005F41 : data <= 8'b00000000 ;
			15'h00005F42 : data <= 8'b00000000 ;
			15'h00005F43 : data <= 8'b00000000 ;
			15'h00005F44 : data <= 8'b00000000 ;
			15'h00005F45 : data <= 8'b00000000 ;
			15'h00005F46 : data <= 8'b00000000 ;
			15'h00005F47 : data <= 8'b00000000 ;
			15'h00005F48 : data <= 8'b00000000 ;
			15'h00005F49 : data <= 8'b00000000 ;
			15'h00005F4A : data <= 8'b00000000 ;
			15'h00005F4B : data <= 8'b00000000 ;
			15'h00005F4C : data <= 8'b00000000 ;
			15'h00005F4D : data <= 8'b00000000 ;
			15'h00005F4E : data <= 8'b00000000 ;
			15'h00005F4F : data <= 8'b00000000 ;
			15'h00005F50 : data <= 8'b00000000 ;
			15'h00005F51 : data <= 8'b00000000 ;
			15'h00005F52 : data <= 8'b00000000 ;
			15'h00005F53 : data <= 8'b00000000 ;
			15'h00005F54 : data <= 8'b00000000 ;
			15'h00005F55 : data <= 8'b00000000 ;
			15'h00005F56 : data <= 8'b00000000 ;
			15'h00005F57 : data <= 8'b00000000 ;
			15'h00005F58 : data <= 8'b00000000 ;
			15'h00005F59 : data <= 8'b00000000 ;
			15'h00005F5A : data <= 8'b00000000 ;
			15'h00005F5B : data <= 8'b00000000 ;
			15'h00005F5C : data <= 8'b00000000 ;
			15'h00005F5D : data <= 8'b00000000 ;
			15'h00005F5E : data <= 8'b00000000 ;
			15'h00005F5F : data <= 8'b00000000 ;
			15'h00005F60 : data <= 8'b00000000 ;
			15'h00005F61 : data <= 8'b00000000 ;
			15'h00005F62 : data <= 8'b00000000 ;
			15'h00005F63 : data <= 8'b00000000 ;
			15'h00005F64 : data <= 8'b00000000 ;
			15'h00005F65 : data <= 8'b00000000 ;
			15'h00005F66 : data <= 8'b00000000 ;
			15'h00005F67 : data <= 8'b00000000 ;
			15'h00005F68 : data <= 8'b00000000 ;
			15'h00005F69 : data <= 8'b00000000 ;
			15'h00005F6A : data <= 8'b00000000 ;
			15'h00005F6B : data <= 8'b00000000 ;
			15'h00005F6C : data <= 8'b00000000 ;
			15'h00005F6D : data <= 8'b00000000 ;
			15'h00005F6E : data <= 8'b00000000 ;
			15'h00005F6F : data <= 8'b00000000 ;
			15'h00005F70 : data <= 8'b00000000 ;
			15'h00005F71 : data <= 8'b00000000 ;
			15'h00005F72 : data <= 8'b00000000 ;
			15'h00005F73 : data <= 8'b00000000 ;
			15'h00005F74 : data <= 8'b00000000 ;
			15'h00005F75 : data <= 8'b00000000 ;
			15'h00005F76 : data <= 8'b00000000 ;
			15'h00005F77 : data <= 8'b00000000 ;
			15'h00005F78 : data <= 8'b00000000 ;
			15'h00005F79 : data <= 8'b00000000 ;
			15'h00005F7A : data <= 8'b00000000 ;
			15'h00005F7B : data <= 8'b00000000 ;
			15'h00005F7C : data <= 8'b00000000 ;
			15'h00005F7D : data <= 8'b00000000 ;
			15'h00005F7E : data <= 8'b00000000 ;
			15'h00005F7F : data <= 8'b00000000 ;
			15'h00005F80 : data <= 8'b00000000 ;
			15'h00005F81 : data <= 8'b00000000 ;
			15'h00005F82 : data <= 8'b00000000 ;
			15'h00005F83 : data <= 8'b00000000 ;
			15'h00005F84 : data <= 8'b00000000 ;
			15'h00005F85 : data <= 8'b00000000 ;
			15'h00005F86 : data <= 8'b00000000 ;
			15'h00005F87 : data <= 8'b00000000 ;
			15'h00005F88 : data <= 8'b00000000 ;
			15'h00005F89 : data <= 8'b00000000 ;
			15'h00005F8A : data <= 8'b00000000 ;
			15'h00005F8B : data <= 8'b00000000 ;
			15'h00005F8C : data <= 8'b00000000 ;
			15'h00005F8D : data <= 8'b00000000 ;
			15'h00005F8E : data <= 8'b00000000 ;
			15'h00005F8F : data <= 8'b00000000 ;
			15'h00005F90 : data <= 8'b00000000 ;
			15'h00005F91 : data <= 8'b00000000 ;
			15'h00005F92 : data <= 8'b00000000 ;
			15'h00005F93 : data <= 8'b00000000 ;
			15'h00005F94 : data <= 8'b00000000 ;
			15'h00005F95 : data <= 8'b00000000 ;
			15'h00005F96 : data <= 8'b00000000 ;
			15'h00005F97 : data <= 8'b00000000 ;
			15'h00005F98 : data <= 8'b00000000 ;
			15'h00005F99 : data <= 8'b00000000 ;
			15'h00005F9A : data <= 8'b00000000 ;
			15'h00005F9B : data <= 8'b00000000 ;
			15'h00005F9C : data <= 8'b00000000 ;
			15'h00005F9D : data <= 8'b00000000 ;
			15'h00005F9E : data <= 8'b00000000 ;
			15'h00005F9F : data <= 8'b00000000 ;
			15'h00005FA0 : data <= 8'b00000000 ;
			15'h00005FA1 : data <= 8'b00000000 ;
			15'h00005FA2 : data <= 8'b00000000 ;
			15'h00005FA3 : data <= 8'b00000000 ;
			15'h00005FA4 : data <= 8'b00000000 ;
			15'h00005FA5 : data <= 8'b00000000 ;
			15'h00005FA6 : data <= 8'b00000000 ;
			15'h00005FA7 : data <= 8'b00000000 ;
			15'h00005FA8 : data <= 8'b00000000 ;
			15'h00005FA9 : data <= 8'b00000000 ;
			15'h00005FAA : data <= 8'b00000000 ;
			15'h00005FAB : data <= 8'b00000000 ;
			15'h00005FAC : data <= 8'b00000000 ;
			15'h00005FAD : data <= 8'b00000000 ;
			15'h00005FAE : data <= 8'b00000000 ;
			15'h00005FAF : data <= 8'b00000000 ;
			15'h00005FB0 : data <= 8'b00000000 ;
			15'h00005FB1 : data <= 8'b00000000 ;
			15'h00005FB2 : data <= 8'b00000000 ;
			15'h00005FB3 : data <= 8'b00000000 ;
			15'h00005FB4 : data <= 8'b00000000 ;
			15'h00005FB5 : data <= 8'b00000000 ;
			15'h00005FB6 : data <= 8'b00000000 ;
			15'h00005FB7 : data <= 8'b00000000 ;
			15'h00005FB8 : data <= 8'b00000000 ;
			15'h00005FB9 : data <= 8'b00000000 ;
			15'h00005FBA : data <= 8'b00000000 ;
			15'h00005FBB : data <= 8'b00000000 ;
			15'h00005FBC : data <= 8'b00000000 ;
			15'h00005FBD : data <= 8'b00000000 ;
			15'h00005FBE : data <= 8'b00000000 ;
			15'h00005FBF : data <= 8'b00000000 ;
			15'h00005FC0 : data <= 8'b00000000 ;
			15'h00005FC1 : data <= 8'b00000000 ;
			15'h00005FC2 : data <= 8'b00000000 ;
			15'h00005FC3 : data <= 8'b00000000 ;
			15'h00005FC4 : data <= 8'b00000000 ;
			15'h00005FC5 : data <= 8'b00000000 ;
			15'h00005FC6 : data <= 8'b00000000 ;
			15'h00005FC7 : data <= 8'b00000000 ;
			15'h00005FC8 : data <= 8'b00000000 ;
			15'h00005FC9 : data <= 8'b00000000 ;
			15'h00005FCA : data <= 8'b00000000 ;
			15'h00005FCB : data <= 8'b00000000 ;
			15'h00005FCC : data <= 8'b00000000 ;
			15'h00005FCD : data <= 8'b00000000 ;
			15'h00005FCE : data <= 8'b00000000 ;
			15'h00005FCF : data <= 8'b00000000 ;
			15'h00005FD0 : data <= 8'b00000000 ;
			15'h00005FD1 : data <= 8'b00000000 ;
			15'h00005FD2 : data <= 8'b00000000 ;
			15'h00005FD3 : data <= 8'b00000000 ;
			15'h00005FD4 : data <= 8'b00000000 ;
			15'h00005FD5 : data <= 8'b00000000 ;
			15'h00005FD6 : data <= 8'b00000000 ;
			15'h00005FD7 : data <= 8'b00000000 ;
			15'h00005FD8 : data <= 8'b00000000 ;
			15'h00005FD9 : data <= 8'b00000000 ;
			15'h00005FDA : data <= 8'b00000000 ;
			15'h00005FDB : data <= 8'b00000000 ;
			15'h00005FDC : data <= 8'b00000000 ;
			15'h00005FDD : data <= 8'b00000000 ;
			15'h00005FDE : data <= 8'b00000000 ;
			15'h00005FDF : data <= 8'b00000000 ;
			15'h00005FE0 : data <= 8'b00000000 ;
			15'h00005FE1 : data <= 8'b00000000 ;
			15'h00005FE2 : data <= 8'b00000000 ;
			15'h00005FE3 : data <= 8'b00000000 ;
			15'h00005FE4 : data <= 8'b00000000 ;
			15'h00005FE5 : data <= 8'b00000000 ;
			15'h00005FE6 : data <= 8'b00000000 ;
			15'h00005FE7 : data <= 8'b00000000 ;
			15'h00005FE8 : data <= 8'b00000000 ;
			15'h00005FE9 : data <= 8'b00000000 ;
			15'h00005FEA : data <= 8'b00000000 ;
			15'h00005FEB : data <= 8'b00000000 ;
			15'h00005FEC : data <= 8'b00000000 ;
			15'h00005FED : data <= 8'b00000000 ;
			15'h00005FEE : data <= 8'b00000000 ;
			15'h00005FEF : data <= 8'b00000000 ;
			15'h00005FF0 : data <= 8'b00000000 ;
			15'h00005FF1 : data <= 8'b00000000 ;
			15'h00005FF2 : data <= 8'b00000000 ;
			15'h00005FF3 : data <= 8'b00000000 ;
			15'h00005FF4 : data <= 8'b00000000 ;
			15'h00005FF5 : data <= 8'b00000000 ;
			15'h00005FF6 : data <= 8'b00000000 ;
			15'h00005FF7 : data <= 8'b00000000 ;
			15'h00005FF8 : data <= 8'b00000000 ;
			15'h00005FF9 : data <= 8'b00000000 ;
			15'h00005FFA : data <= 8'b00000000 ;
			15'h00005FFB : data <= 8'b00000000 ;
			15'h00005FFC : data <= 8'b00000000 ;
			15'h00005FFD : data <= 8'b00000000 ;
			15'h00005FFE : data <= 8'b00000000 ;
			15'h00005FFF : data <= 8'b00000000 ;
			15'h00006000 : data <= 8'b00000000 ;
			15'h00006001 : data <= 8'b00000000 ;
			15'h00006002 : data <= 8'b00000000 ;
			15'h00006003 : data <= 8'b00000000 ;
			15'h00006004 : data <= 8'b00000000 ;
			15'h00006005 : data <= 8'b00000000 ;
			15'h00006006 : data <= 8'b00000000 ;
			15'h00006007 : data <= 8'b00000000 ;
			15'h00006008 : data <= 8'b00000000 ;
			15'h00006009 : data <= 8'b00000000 ;
			15'h0000600A : data <= 8'b00000000 ;
			15'h0000600B : data <= 8'b00000000 ;
			15'h0000600C : data <= 8'b00000000 ;
			15'h0000600D : data <= 8'b00000000 ;
			15'h0000600E : data <= 8'b00000000 ;
			15'h0000600F : data <= 8'b00000000 ;
			15'h00006010 : data <= 8'b00000000 ;
			15'h00006011 : data <= 8'b00000000 ;
			15'h00006012 : data <= 8'b00000000 ;
			15'h00006013 : data <= 8'b00000000 ;
			15'h00006014 : data <= 8'b00000000 ;
			15'h00006015 : data <= 8'b00000000 ;
			15'h00006016 : data <= 8'b00000000 ;
			15'h00006017 : data <= 8'b00000000 ;
			15'h00006018 : data <= 8'b00000000 ;
			15'h00006019 : data <= 8'b00000000 ;
			15'h0000601A : data <= 8'b00000000 ;
			15'h0000601B : data <= 8'b00000000 ;
			15'h0000601C : data <= 8'b00000000 ;
			15'h0000601D : data <= 8'b00000000 ;
			15'h0000601E : data <= 8'b00000000 ;
			15'h0000601F : data <= 8'b00000000 ;
			15'h00006020 : data <= 8'b00000000 ;
			15'h00006021 : data <= 8'b00000000 ;
			15'h00006022 : data <= 8'b00000000 ;
			15'h00006023 : data <= 8'b00000000 ;
			15'h00006024 : data <= 8'b00000000 ;
			15'h00006025 : data <= 8'b00000000 ;
			15'h00006026 : data <= 8'b00000000 ;
			15'h00006027 : data <= 8'b00000000 ;
			15'h00006028 : data <= 8'b00000000 ;
			15'h00006029 : data <= 8'b00000000 ;
			15'h0000602A : data <= 8'b00000000 ;
			15'h0000602B : data <= 8'b00000000 ;
			15'h0000602C : data <= 8'b00000000 ;
			15'h0000602D : data <= 8'b00000000 ;
			15'h0000602E : data <= 8'b00000000 ;
			15'h0000602F : data <= 8'b00000000 ;
			15'h00006030 : data <= 8'b00000000 ;
			15'h00006031 : data <= 8'b00000000 ;
			15'h00006032 : data <= 8'b00000000 ;
			15'h00006033 : data <= 8'b00000000 ;
			15'h00006034 : data <= 8'b00000000 ;
			15'h00006035 : data <= 8'b00000000 ;
			15'h00006036 : data <= 8'b00000000 ;
			15'h00006037 : data <= 8'b00000000 ;
			15'h00006038 : data <= 8'b00000000 ;
			15'h00006039 : data <= 8'b00000000 ;
			15'h0000603A : data <= 8'b00000000 ;
			15'h0000603B : data <= 8'b00000000 ;
			15'h0000603C : data <= 8'b00000000 ;
			15'h0000603D : data <= 8'b00000000 ;
			15'h0000603E : data <= 8'b00000000 ;
			15'h0000603F : data <= 8'b00000000 ;
			15'h00006040 : data <= 8'b00000000 ;
			15'h00006041 : data <= 8'b00000000 ;
			15'h00006042 : data <= 8'b00000000 ;
			15'h00006043 : data <= 8'b00000000 ;
			15'h00006044 : data <= 8'b00000000 ;
			15'h00006045 : data <= 8'b00000000 ;
			15'h00006046 : data <= 8'b00000000 ;
			15'h00006047 : data <= 8'b00000000 ;
			15'h00006048 : data <= 8'b00000000 ;
			15'h00006049 : data <= 8'b00000000 ;
			15'h0000604A : data <= 8'b00000000 ;
			15'h0000604B : data <= 8'b00000000 ;
			15'h0000604C : data <= 8'b00000000 ;
			15'h0000604D : data <= 8'b00000000 ;
			15'h0000604E : data <= 8'b00000000 ;
			15'h0000604F : data <= 8'b00000000 ;
			15'h00006050 : data <= 8'b00000000 ;
			15'h00006051 : data <= 8'b00000000 ;
			15'h00006052 : data <= 8'b00000000 ;
			15'h00006053 : data <= 8'b00000000 ;
			15'h00006054 : data <= 8'b00000000 ;
			15'h00006055 : data <= 8'b00000000 ;
			15'h00006056 : data <= 8'b00000000 ;
			15'h00006057 : data <= 8'b00000000 ;
			15'h00006058 : data <= 8'b00000000 ;
			15'h00006059 : data <= 8'b00000000 ;
			15'h0000605A : data <= 8'b00000000 ;
			15'h0000605B : data <= 8'b00000000 ;
			15'h0000605C : data <= 8'b00000000 ;
			15'h0000605D : data <= 8'b00000000 ;
			15'h0000605E : data <= 8'b00000000 ;
			15'h0000605F : data <= 8'b00000000 ;
			15'h00006060 : data <= 8'b00000000 ;
			15'h00006061 : data <= 8'b00000000 ;
			15'h00006062 : data <= 8'b00000000 ;
			15'h00006063 : data <= 8'b00000000 ;
			15'h00006064 : data <= 8'b00000000 ;
			15'h00006065 : data <= 8'b00000000 ;
			15'h00006066 : data <= 8'b00000000 ;
			15'h00006067 : data <= 8'b00000000 ;
			15'h00006068 : data <= 8'b00000000 ;
			15'h00006069 : data <= 8'b00000000 ;
			15'h0000606A : data <= 8'b00000000 ;
			15'h0000606B : data <= 8'b00000000 ;
			15'h0000606C : data <= 8'b00000000 ;
			15'h0000606D : data <= 8'b00000000 ;
			15'h0000606E : data <= 8'b00000000 ;
			15'h0000606F : data <= 8'b00000000 ;
			15'h00006070 : data <= 8'b00000000 ;
			15'h00006071 : data <= 8'b00000000 ;
			15'h00006072 : data <= 8'b00000000 ;
			15'h00006073 : data <= 8'b00000000 ;
			15'h00006074 : data <= 8'b00000000 ;
			15'h00006075 : data <= 8'b00000000 ;
			15'h00006076 : data <= 8'b00000000 ;
			15'h00006077 : data <= 8'b00000000 ;
			15'h00006078 : data <= 8'b00000000 ;
			15'h00006079 : data <= 8'b00000000 ;
			15'h0000607A : data <= 8'b00000000 ;
			15'h0000607B : data <= 8'b00000000 ;
			15'h0000607C : data <= 8'b00000000 ;
			15'h0000607D : data <= 8'b00000000 ;
			15'h0000607E : data <= 8'b00000000 ;
			15'h0000607F : data <= 8'b00000000 ;
			15'h00006080 : data <= 8'b00000000 ;
			15'h00006081 : data <= 8'b00000000 ;
			15'h00006082 : data <= 8'b00000000 ;
			15'h00006083 : data <= 8'b00000000 ;
			15'h00006084 : data <= 8'b00000000 ;
			15'h00006085 : data <= 8'b00000000 ;
			15'h00006086 : data <= 8'b00000000 ;
			15'h00006087 : data <= 8'b00000000 ;
			15'h00006088 : data <= 8'b00000000 ;
			15'h00006089 : data <= 8'b00000000 ;
			15'h0000608A : data <= 8'b00000000 ;
			15'h0000608B : data <= 8'b00000000 ;
			15'h0000608C : data <= 8'b00000000 ;
			15'h0000608D : data <= 8'b00000000 ;
			15'h0000608E : data <= 8'b00000000 ;
			15'h0000608F : data <= 8'b00000000 ;
			15'h00006090 : data <= 8'b00000000 ;
			15'h00006091 : data <= 8'b00000000 ;
			15'h00006092 : data <= 8'b00000000 ;
			15'h00006093 : data <= 8'b00000000 ;
			15'h00006094 : data <= 8'b00000000 ;
			15'h00006095 : data <= 8'b00000000 ;
			15'h00006096 : data <= 8'b00000000 ;
			15'h00006097 : data <= 8'b00000000 ;
			15'h00006098 : data <= 8'b00000000 ;
			15'h00006099 : data <= 8'b00000000 ;
			15'h0000609A : data <= 8'b00000000 ;
			15'h0000609B : data <= 8'b00000000 ;
			15'h0000609C : data <= 8'b00000000 ;
			15'h0000609D : data <= 8'b00000000 ;
			15'h0000609E : data <= 8'b00000000 ;
			15'h0000609F : data <= 8'b00000000 ;
			15'h000060A0 : data <= 8'b00000000 ;
			15'h000060A1 : data <= 8'b00000000 ;
			15'h000060A2 : data <= 8'b00000000 ;
			15'h000060A3 : data <= 8'b00000000 ;
			15'h000060A4 : data <= 8'b00000000 ;
			15'h000060A5 : data <= 8'b00000000 ;
			15'h000060A6 : data <= 8'b00000000 ;
			15'h000060A7 : data <= 8'b00000000 ;
			15'h000060A8 : data <= 8'b00000000 ;
			15'h000060A9 : data <= 8'b00000000 ;
			15'h000060AA : data <= 8'b00000000 ;
			15'h000060AB : data <= 8'b00000000 ;
			15'h000060AC : data <= 8'b00000000 ;
			15'h000060AD : data <= 8'b00000000 ;
			15'h000060AE : data <= 8'b00000000 ;
			15'h000060AF : data <= 8'b00000000 ;
			15'h000060B0 : data <= 8'b00000000 ;
			15'h000060B1 : data <= 8'b00000000 ;
			15'h000060B2 : data <= 8'b00000000 ;
			15'h000060B3 : data <= 8'b00000000 ;
			15'h000060B4 : data <= 8'b00000000 ;
			15'h000060B5 : data <= 8'b00000000 ;
			15'h000060B6 : data <= 8'b00000000 ;
			15'h000060B7 : data <= 8'b00000000 ;
			15'h000060B8 : data <= 8'b00000000 ;
			15'h000060B9 : data <= 8'b00000000 ;
			15'h000060BA : data <= 8'b00000000 ;
			15'h000060BB : data <= 8'b00000000 ;
			15'h000060BC : data <= 8'b00000000 ;
			15'h000060BD : data <= 8'b00000000 ;
			15'h000060BE : data <= 8'b00000000 ;
			15'h000060BF : data <= 8'b00000000 ;
			15'h000060C0 : data <= 8'b00000000 ;
			15'h000060C1 : data <= 8'b00000000 ;
			15'h000060C2 : data <= 8'b00000000 ;
			15'h000060C3 : data <= 8'b00000000 ;
			15'h000060C4 : data <= 8'b00000000 ;
			15'h000060C5 : data <= 8'b00000000 ;
			15'h000060C6 : data <= 8'b00000000 ;
			15'h000060C7 : data <= 8'b00000000 ;
			15'h000060C8 : data <= 8'b00000000 ;
			15'h000060C9 : data <= 8'b00000000 ;
			15'h000060CA : data <= 8'b00000000 ;
			15'h000060CB : data <= 8'b00000000 ;
			15'h000060CC : data <= 8'b00000000 ;
			15'h000060CD : data <= 8'b00000000 ;
			15'h000060CE : data <= 8'b00000000 ;
			15'h000060CF : data <= 8'b00000000 ;
			15'h000060D0 : data <= 8'b00000000 ;
			15'h000060D1 : data <= 8'b00000000 ;
			15'h000060D2 : data <= 8'b00000000 ;
			15'h000060D3 : data <= 8'b00000000 ;
			15'h000060D4 : data <= 8'b00000000 ;
			15'h000060D5 : data <= 8'b00000000 ;
			15'h000060D6 : data <= 8'b00000000 ;
			15'h000060D7 : data <= 8'b00000000 ;
			15'h000060D8 : data <= 8'b00000000 ;
			15'h000060D9 : data <= 8'b00000000 ;
			15'h000060DA : data <= 8'b00000000 ;
			15'h000060DB : data <= 8'b00000000 ;
			15'h000060DC : data <= 8'b00000000 ;
			15'h000060DD : data <= 8'b00000000 ;
			15'h000060DE : data <= 8'b00000000 ;
			15'h000060DF : data <= 8'b00000000 ;
			15'h000060E0 : data <= 8'b00000000 ;
			15'h000060E1 : data <= 8'b00000000 ;
			15'h000060E2 : data <= 8'b00000000 ;
			15'h000060E3 : data <= 8'b00000000 ;
			15'h000060E4 : data <= 8'b00000000 ;
			15'h000060E5 : data <= 8'b00000000 ;
			15'h000060E6 : data <= 8'b00000000 ;
			15'h000060E7 : data <= 8'b00000000 ;
			15'h000060E8 : data <= 8'b00000000 ;
			15'h000060E9 : data <= 8'b00000000 ;
			15'h000060EA : data <= 8'b00000000 ;
			15'h000060EB : data <= 8'b00000000 ;
			15'h000060EC : data <= 8'b00000000 ;
			15'h000060ED : data <= 8'b00000000 ;
			15'h000060EE : data <= 8'b00000000 ;
			15'h000060EF : data <= 8'b00000000 ;
			15'h000060F0 : data <= 8'b00000000 ;
			15'h000060F1 : data <= 8'b00000000 ;
			15'h000060F2 : data <= 8'b00000000 ;
			15'h000060F3 : data <= 8'b00000000 ;
			15'h000060F4 : data <= 8'b00000000 ;
			15'h000060F5 : data <= 8'b00000000 ;
			15'h000060F6 : data <= 8'b00000000 ;
			15'h000060F7 : data <= 8'b00000000 ;
			15'h000060F8 : data <= 8'b00000000 ;
			15'h000060F9 : data <= 8'b00000000 ;
			15'h000060FA : data <= 8'b00000000 ;
			15'h000060FB : data <= 8'b00000000 ;
			15'h000060FC : data <= 8'b00000000 ;
			15'h000060FD : data <= 8'b00000000 ;
			15'h000060FE : data <= 8'b00000000 ;
			15'h000060FF : data <= 8'b00000000 ;
			15'h00006100 : data <= 8'b00000000 ;
			15'h00006101 : data <= 8'b00000000 ;
			15'h00006102 : data <= 8'b00000000 ;
			15'h00006103 : data <= 8'b00000000 ;
			15'h00006104 : data <= 8'b00000000 ;
			15'h00006105 : data <= 8'b00000000 ;
			15'h00006106 : data <= 8'b00000000 ;
			15'h00006107 : data <= 8'b00000000 ;
			15'h00006108 : data <= 8'b00000000 ;
			15'h00006109 : data <= 8'b00000000 ;
			15'h0000610A : data <= 8'b00000000 ;
			15'h0000610B : data <= 8'b00000000 ;
			15'h0000610C : data <= 8'b00000000 ;
			15'h0000610D : data <= 8'b00000000 ;
			15'h0000610E : data <= 8'b00000000 ;
			15'h0000610F : data <= 8'b00000000 ;
			15'h00006110 : data <= 8'b00000000 ;
			15'h00006111 : data <= 8'b00000000 ;
			15'h00006112 : data <= 8'b00000000 ;
			15'h00006113 : data <= 8'b00000000 ;
			15'h00006114 : data <= 8'b00000000 ;
			15'h00006115 : data <= 8'b00000000 ;
			15'h00006116 : data <= 8'b00000000 ;
			15'h00006117 : data <= 8'b00000000 ;
			15'h00006118 : data <= 8'b00000000 ;
			15'h00006119 : data <= 8'b00000000 ;
			15'h0000611A : data <= 8'b00000000 ;
			15'h0000611B : data <= 8'b00000000 ;
			15'h0000611C : data <= 8'b00000000 ;
			15'h0000611D : data <= 8'b00000000 ;
			15'h0000611E : data <= 8'b00000000 ;
			15'h0000611F : data <= 8'b00000000 ;
			15'h00006120 : data <= 8'b00000000 ;
			15'h00006121 : data <= 8'b00000000 ;
			15'h00006122 : data <= 8'b00000000 ;
			15'h00006123 : data <= 8'b00000000 ;
			15'h00006124 : data <= 8'b00000000 ;
			15'h00006125 : data <= 8'b00000000 ;
			15'h00006126 : data <= 8'b00000000 ;
			15'h00006127 : data <= 8'b00000000 ;
			15'h00006128 : data <= 8'b00000000 ;
			15'h00006129 : data <= 8'b00000000 ;
			15'h0000612A : data <= 8'b00000000 ;
			15'h0000612B : data <= 8'b00000000 ;
			15'h0000612C : data <= 8'b00000000 ;
			15'h0000612D : data <= 8'b00000000 ;
			15'h0000612E : data <= 8'b00000000 ;
			15'h0000612F : data <= 8'b00000000 ;
			15'h00006130 : data <= 8'b00000000 ;
			15'h00006131 : data <= 8'b00000000 ;
			15'h00006132 : data <= 8'b00000000 ;
			15'h00006133 : data <= 8'b00000000 ;
			15'h00006134 : data <= 8'b00000000 ;
			15'h00006135 : data <= 8'b00000000 ;
			15'h00006136 : data <= 8'b00000000 ;
			15'h00006137 : data <= 8'b00000000 ;
			15'h00006138 : data <= 8'b00000000 ;
			15'h00006139 : data <= 8'b00000000 ;
			15'h0000613A : data <= 8'b00000000 ;
			15'h0000613B : data <= 8'b00000000 ;
			15'h0000613C : data <= 8'b00000000 ;
			15'h0000613D : data <= 8'b00000000 ;
			15'h0000613E : data <= 8'b00000000 ;
			15'h0000613F : data <= 8'b00000000 ;
			15'h00006140 : data <= 8'b00000000 ;
			15'h00006141 : data <= 8'b00000000 ;
			15'h00006142 : data <= 8'b00000000 ;
			15'h00006143 : data <= 8'b00000000 ;
			15'h00006144 : data <= 8'b00000000 ;
			15'h00006145 : data <= 8'b00000000 ;
			15'h00006146 : data <= 8'b00000000 ;
			15'h00006147 : data <= 8'b00000000 ;
			15'h00006148 : data <= 8'b00000000 ;
			15'h00006149 : data <= 8'b00000000 ;
			15'h0000614A : data <= 8'b00000000 ;
			15'h0000614B : data <= 8'b00000000 ;
			15'h0000614C : data <= 8'b00000000 ;
			15'h0000614D : data <= 8'b00000000 ;
			15'h0000614E : data <= 8'b00000000 ;
			15'h0000614F : data <= 8'b00000000 ;
			15'h00006150 : data <= 8'b00000000 ;
			15'h00006151 : data <= 8'b00000000 ;
			15'h00006152 : data <= 8'b00000000 ;
			15'h00006153 : data <= 8'b00000000 ;
			15'h00006154 : data <= 8'b00000000 ;
			15'h00006155 : data <= 8'b00000000 ;
			15'h00006156 : data <= 8'b00000000 ;
			15'h00006157 : data <= 8'b00000000 ;
			15'h00006158 : data <= 8'b00000000 ;
			15'h00006159 : data <= 8'b00000000 ;
			15'h0000615A : data <= 8'b00000000 ;
			15'h0000615B : data <= 8'b00000000 ;
			15'h0000615C : data <= 8'b00000000 ;
			15'h0000615D : data <= 8'b00000000 ;
			15'h0000615E : data <= 8'b00000000 ;
			15'h0000615F : data <= 8'b00000000 ;
			15'h00006160 : data <= 8'b00000000 ;
			15'h00006161 : data <= 8'b00000000 ;
			15'h00006162 : data <= 8'b00000000 ;
			15'h00006163 : data <= 8'b00000000 ;
			15'h00006164 : data <= 8'b00000000 ;
			15'h00006165 : data <= 8'b00000000 ;
			15'h00006166 : data <= 8'b00000000 ;
			15'h00006167 : data <= 8'b00000000 ;
			15'h00006168 : data <= 8'b00000000 ;
			15'h00006169 : data <= 8'b00000000 ;
			15'h0000616A : data <= 8'b00000000 ;
			15'h0000616B : data <= 8'b00000000 ;
			15'h0000616C : data <= 8'b00000000 ;
			15'h0000616D : data <= 8'b00000000 ;
			15'h0000616E : data <= 8'b00000000 ;
			15'h0000616F : data <= 8'b00000000 ;
			15'h00006170 : data <= 8'b00000000 ;
			15'h00006171 : data <= 8'b00000000 ;
			15'h00006172 : data <= 8'b00000000 ;
			15'h00006173 : data <= 8'b00000000 ;
			15'h00006174 : data <= 8'b00000000 ;
			15'h00006175 : data <= 8'b00000000 ;
			15'h00006176 : data <= 8'b00000000 ;
			15'h00006177 : data <= 8'b00000000 ;
			15'h00006178 : data <= 8'b00000000 ;
			15'h00006179 : data <= 8'b00000000 ;
			15'h0000617A : data <= 8'b00000000 ;
			15'h0000617B : data <= 8'b00000000 ;
			15'h0000617C : data <= 8'b00000000 ;
			15'h0000617D : data <= 8'b00000000 ;
			15'h0000617E : data <= 8'b00000000 ;
			15'h0000617F : data <= 8'b00000000 ;
			15'h00006180 : data <= 8'b00000000 ;
			15'h00006181 : data <= 8'b00000000 ;
			15'h00006182 : data <= 8'b00000000 ;
			15'h00006183 : data <= 8'b00000000 ;
			15'h00006184 : data <= 8'b00000000 ;
			15'h00006185 : data <= 8'b00000000 ;
			15'h00006186 : data <= 8'b00000000 ;
			15'h00006187 : data <= 8'b00000000 ;
			15'h00006188 : data <= 8'b00000000 ;
			15'h00006189 : data <= 8'b00000000 ;
			15'h0000618A : data <= 8'b00000000 ;
			15'h0000618B : data <= 8'b00000000 ;
			15'h0000618C : data <= 8'b00000000 ;
			15'h0000618D : data <= 8'b00000000 ;
			15'h0000618E : data <= 8'b00000000 ;
			15'h0000618F : data <= 8'b00000000 ;
			15'h00006190 : data <= 8'b00000000 ;
			15'h00006191 : data <= 8'b00000000 ;
			15'h00006192 : data <= 8'b00000000 ;
			15'h00006193 : data <= 8'b00000000 ;
			15'h00006194 : data <= 8'b00000000 ;
			15'h00006195 : data <= 8'b00000000 ;
			15'h00006196 : data <= 8'b00000000 ;
			15'h00006197 : data <= 8'b00000000 ;
			15'h00006198 : data <= 8'b00000000 ;
			15'h00006199 : data <= 8'b00000000 ;
			15'h0000619A : data <= 8'b00000000 ;
			15'h0000619B : data <= 8'b00000000 ;
			15'h0000619C : data <= 8'b00000000 ;
			15'h0000619D : data <= 8'b00000000 ;
			15'h0000619E : data <= 8'b00000000 ;
			15'h0000619F : data <= 8'b00000000 ;
			15'h000061A0 : data <= 8'b00000000 ;
			15'h000061A1 : data <= 8'b00000000 ;
			15'h000061A2 : data <= 8'b00000000 ;
			15'h000061A3 : data <= 8'b00000000 ;
			15'h000061A4 : data <= 8'b00000000 ;
			15'h000061A5 : data <= 8'b00000000 ;
			15'h000061A6 : data <= 8'b00000000 ;
			15'h000061A7 : data <= 8'b00000000 ;
			15'h000061A8 : data <= 8'b00000000 ;
			15'h000061A9 : data <= 8'b00000000 ;
			15'h000061AA : data <= 8'b00000000 ;
			15'h000061AB : data <= 8'b00000000 ;
			15'h000061AC : data <= 8'b00000000 ;
			15'h000061AD : data <= 8'b00000000 ;
			15'h000061AE : data <= 8'b00000000 ;
			15'h000061AF : data <= 8'b00000000 ;
			15'h000061B0 : data <= 8'b00000000 ;
			15'h000061B1 : data <= 8'b00000000 ;
			15'h000061B2 : data <= 8'b00000000 ;
			15'h000061B3 : data <= 8'b00000000 ;
			15'h000061B4 : data <= 8'b00000000 ;
			15'h000061B5 : data <= 8'b00000000 ;
			15'h000061B6 : data <= 8'b00000000 ;
			15'h000061B7 : data <= 8'b00000000 ;
			15'h000061B8 : data <= 8'b00000000 ;
			15'h000061B9 : data <= 8'b00000000 ;
			15'h000061BA : data <= 8'b00000000 ;
			15'h000061BB : data <= 8'b00000000 ;
			15'h000061BC : data <= 8'b00000000 ;
			15'h000061BD : data <= 8'b00000000 ;
			15'h000061BE : data <= 8'b00000000 ;
			15'h000061BF : data <= 8'b00000000 ;
			15'h000061C0 : data <= 8'b00000000 ;
			15'h000061C1 : data <= 8'b00000000 ;
			15'h000061C2 : data <= 8'b00000000 ;
			15'h000061C3 : data <= 8'b00000000 ;
			15'h000061C4 : data <= 8'b00000000 ;
			15'h000061C5 : data <= 8'b00000000 ;
			15'h000061C6 : data <= 8'b00000000 ;
			15'h000061C7 : data <= 8'b00000000 ;
			15'h000061C8 : data <= 8'b00000000 ;
			15'h000061C9 : data <= 8'b00000000 ;
			15'h000061CA : data <= 8'b00000000 ;
			15'h000061CB : data <= 8'b00000000 ;
			15'h000061CC : data <= 8'b00000000 ;
			15'h000061CD : data <= 8'b00000000 ;
			15'h000061CE : data <= 8'b00000000 ;
			15'h000061CF : data <= 8'b00000000 ;
			15'h000061D0 : data <= 8'b00000000 ;
			15'h000061D1 : data <= 8'b00000000 ;
			15'h000061D2 : data <= 8'b00000000 ;
			15'h000061D3 : data <= 8'b00000000 ;
			15'h000061D4 : data <= 8'b00000000 ;
			15'h000061D5 : data <= 8'b00000000 ;
			15'h000061D6 : data <= 8'b00000000 ;
			15'h000061D7 : data <= 8'b00000000 ;
			15'h000061D8 : data <= 8'b00000000 ;
			15'h000061D9 : data <= 8'b00000000 ;
			15'h000061DA : data <= 8'b00000000 ;
			15'h000061DB : data <= 8'b00000000 ;
			15'h000061DC : data <= 8'b00000000 ;
			15'h000061DD : data <= 8'b00000000 ;
			15'h000061DE : data <= 8'b00000000 ;
			15'h000061DF : data <= 8'b00000000 ;
			15'h000061E0 : data <= 8'b00000000 ;
			15'h000061E1 : data <= 8'b00000000 ;
			15'h000061E2 : data <= 8'b00000000 ;
			15'h000061E3 : data <= 8'b00000000 ;
			15'h000061E4 : data <= 8'b00000000 ;
			15'h000061E5 : data <= 8'b00000000 ;
			15'h000061E6 : data <= 8'b00000000 ;
			15'h000061E7 : data <= 8'b00000000 ;
			15'h000061E8 : data <= 8'b00000000 ;
			15'h000061E9 : data <= 8'b00000000 ;
			15'h000061EA : data <= 8'b00000000 ;
			15'h000061EB : data <= 8'b00000000 ;
			15'h000061EC : data <= 8'b00000000 ;
			15'h000061ED : data <= 8'b00000000 ;
			15'h000061EE : data <= 8'b00000000 ;
			15'h000061EF : data <= 8'b00000000 ;
			15'h000061F0 : data <= 8'b00000000 ;
			15'h000061F1 : data <= 8'b00000000 ;
			15'h000061F2 : data <= 8'b00000000 ;
			15'h000061F3 : data <= 8'b00000000 ;
			15'h000061F4 : data <= 8'b00000000 ;
			15'h000061F5 : data <= 8'b00000000 ;
			15'h000061F6 : data <= 8'b00000000 ;
			15'h000061F7 : data <= 8'b00000000 ;
			15'h000061F8 : data <= 8'b00000000 ;
			15'h000061F9 : data <= 8'b00000000 ;
			15'h000061FA : data <= 8'b00000000 ;
			15'h000061FB : data <= 8'b00000000 ;
			15'h000061FC : data <= 8'b00000000 ;
			15'h000061FD : data <= 8'b00000000 ;
			15'h000061FE : data <= 8'b00000000 ;
			15'h000061FF : data <= 8'b00000000 ;
			15'h00006200 : data <= 8'b00000000 ;
			15'h00006201 : data <= 8'b00000000 ;
			15'h00006202 : data <= 8'b00000000 ;
			15'h00006203 : data <= 8'b00000000 ;
			15'h00006204 : data <= 8'b00000000 ;
			15'h00006205 : data <= 8'b00000000 ;
			15'h00006206 : data <= 8'b00000000 ;
			15'h00006207 : data <= 8'b00000000 ;
			15'h00006208 : data <= 8'b00000000 ;
			15'h00006209 : data <= 8'b00000000 ;
			15'h0000620A : data <= 8'b00000000 ;
			15'h0000620B : data <= 8'b00000000 ;
			15'h0000620C : data <= 8'b00000000 ;
			15'h0000620D : data <= 8'b00000000 ;
			15'h0000620E : data <= 8'b00000000 ;
			15'h0000620F : data <= 8'b00000000 ;
			15'h00006210 : data <= 8'b00000000 ;
			15'h00006211 : data <= 8'b00000000 ;
			15'h00006212 : data <= 8'b00000000 ;
			15'h00006213 : data <= 8'b00000000 ;
			15'h00006214 : data <= 8'b00000000 ;
			15'h00006215 : data <= 8'b00000000 ;
			15'h00006216 : data <= 8'b00000000 ;
			15'h00006217 : data <= 8'b00000000 ;
			15'h00006218 : data <= 8'b00000000 ;
			15'h00006219 : data <= 8'b00000000 ;
			15'h0000621A : data <= 8'b00000000 ;
			15'h0000621B : data <= 8'b00000000 ;
			15'h0000621C : data <= 8'b00000000 ;
			15'h0000621D : data <= 8'b00000000 ;
			15'h0000621E : data <= 8'b00000000 ;
			15'h0000621F : data <= 8'b00000000 ;
			15'h00006220 : data <= 8'b00000000 ;
			15'h00006221 : data <= 8'b00000000 ;
			15'h00006222 : data <= 8'b00000000 ;
			15'h00006223 : data <= 8'b00000000 ;
			15'h00006224 : data <= 8'b00000000 ;
			15'h00006225 : data <= 8'b00000000 ;
			15'h00006226 : data <= 8'b00000000 ;
			15'h00006227 : data <= 8'b00000000 ;
			15'h00006228 : data <= 8'b00000000 ;
			15'h00006229 : data <= 8'b00000000 ;
			15'h0000622A : data <= 8'b00000000 ;
			15'h0000622B : data <= 8'b00000000 ;
			15'h0000622C : data <= 8'b00000000 ;
			15'h0000622D : data <= 8'b00000000 ;
			15'h0000622E : data <= 8'b00000000 ;
			15'h0000622F : data <= 8'b00000000 ;
			15'h00006230 : data <= 8'b00000000 ;
			15'h00006231 : data <= 8'b00000000 ;
			15'h00006232 : data <= 8'b00000000 ;
			15'h00006233 : data <= 8'b00000000 ;
			15'h00006234 : data <= 8'b00000000 ;
			15'h00006235 : data <= 8'b00000000 ;
			15'h00006236 : data <= 8'b00000000 ;
			15'h00006237 : data <= 8'b00000000 ;
			15'h00006238 : data <= 8'b00000000 ;
			15'h00006239 : data <= 8'b00000000 ;
			15'h0000623A : data <= 8'b00000000 ;
			15'h0000623B : data <= 8'b00000000 ;
			15'h0000623C : data <= 8'b00000000 ;
			15'h0000623D : data <= 8'b00000000 ;
			15'h0000623E : data <= 8'b00000000 ;
			15'h0000623F : data <= 8'b00000000 ;
			15'h00006240 : data <= 8'b00000000 ;
			15'h00006241 : data <= 8'b00000000 ;
			15'h00006242 : data <= 8'b00000000 ;
			15'h00006243 : data <= 8'b00000000 ;
			15'h00006244 : data <= 8'b00000000 ;
			15'h00006245 : data <= 8'b00000000 ;
			15'h00006246 : data <= 8'b00000000 ;
			15'h00006247 : data <= 8'b00000000 ;
			15'h00006248 : data <= 8'b00000000 ;
			15'h00006249 : data <= 8'b00000000 ;
			15'h0000624A : data <= 8'b00000000 ;
			15'h0000624B : data <= 8'b00000000 ;
			15'h0000624C : data <= 8'b00000000 ;
			15'h0000624D : data <= 8'b00000000 ;
			15'h0000624E : data <= 8'b00000000 ;
			15'h0000624F : data <= 8'b00000000 ;
			15'h00006250 : data <= 8'b00000000 ;
			15'h00006251 : data <= 8'b00000000 ;
			15'h00006252 : data <= 8'b00000000 ;
			15'h00006253 : data <= 8'b00000000 ;
			15'h00006254 : data <= 8'b00000000 ;
			15'h00006255 : data <= 8'b00000000 ;
			15'h00006256 : data <= 8'b00000000 ;
			15'h00006257 : data <= 8'b00000000 ;
			15'h00006258 : data <= 8'b00000000 ;
			15'h00006259 : data <= 8'b00000000 ;
			15'h0000625A : data <= 8'b00000000 ;
			15'h0000625B : data <= 8'b00000000 ;
			15'h0000625C : data <= 8'b00000000 ;
			15'h0000625D : data <= 8'b00000000 ;
			15'h0000625E : data <= 8'b00000000 ;
			15'h0000625F : data <= 8'b00000000 ;
			15'h00006260 : data <= 8'b00000000 ;
			15'h00006261 : data <= 8'b00000000 ;
			15'h00006262 : data <= 8'b00000000 ;
			15'h00006263 : data <= 8'b00000000 ;
			15'h00006264 : data <= 8'b00000000 ;
			15'h00006265 : data <= 8'b00000000 ;
			15'h00006266 : data <= 8'b00000000 ;
			15'h00006267 : data <= 8'b00000000 ;
			15'h00006268 : data <= 8'b00000000 ;
			15'h00006269 : data <= 8'b00000000 ;
			15'h0000626A : data <= 8'b00000000 ;
			15'h0000626B : data <= 8'b00000000 ;
			15'h0000626C : data <= 8'b00000000 ;
			15'h0000626D : data <= 8'b00000000 ;
			15'h0000626E : data <= 8'b00000000 ;
			15'h0000626F : data <= 8'b00000000 ;
			15'h00006270 : data <= 8'b00000000 ;
			15'h00006271 : data <= 8'b00000000 ;
			15'h00006272 : data <= 8'b00000000 ;
			15'h00006273 : data <= 8'b00000000 ;
			15'h00006274 : data <= 8'b00000000 ;
			15'h00006275 : data <= 8'b00000000 ;
			15'h00006276 : data <= 8'b00000000 ;
			15'h00006277 : data <= 8'b00000000 ;
			15'h00006278 : data <= 8'b00000000 ;
			15'h00006279 : data <= 8'b00000000 ;
			15'h0000627A : data <= 8'b00000000 ;
			15'h0000627B : data <= 8'b00000000 ;
			15'h0000627C : data <= 8'b00000000 ;
			15'h0000627D : data <= 8'b00000000 ;
			15'h0000627E : data <= 8'b00000000 ;
			15'h0000627F : data <= 8'b00000000 ;
			15'h00006280 : data <= 8'b00000000 ;
			15'h00006281 : data <= 8'b00000000 ;
			15'h00006282 : data <= 8'b00000000 ;
			15'h00006283 : data <= 8'b00000000 ;
			15'h00006284 : data <= 8'b00000000 ;
			15'h00006285 : data <= 8'b00000000 ;
			15'h00006286 : data <= 8'b00000000 ;
			15'h00006287 : data <= 8'b00000000 ;
			15'h00006288 : data <= 8'b00000000 ;
			15'h00006289 : data <= 8'b00000000 ;
			15'h0000628A : data <= 8'b00000000 ;
			15'h0000628B : data <= 8'b00000000 ;
			15'h0000628C : data <= 8'b00000000 ;
			15'h0000628D : data <= 8'b00000000 ;
			15'h0000628E : data <= 8'b00000000 ;
			15'h0000628F : data <= 8'b00000000 ;
			15'h00006290 : data <= 8'b00000000 ;
			15'h00006291 : data <= 8'b00000000 ;
			15'h00006292 : data <= 8'b00000000 ;
			15'h00006293 : data <= 8'b00000000 ;
			15'h00006294 : data <= 8'b00000000 ;
			15'h00006295 : data <= 8'b00000000 ;
			15'h00006296 : data <= 8'b00000000 ;
			15'h00006297 : data <= 8'b00000000 ;
			15'h00006298 : data <= 8'b00000000 ;
			15'h00006299 : data <= 8'b00000000 ;
			15'h0000629A : data <= 8'b00000000 ;
			15'h0000629B : data <= 8'b00000000 ;
			15'h0000629C : data <= 8'b00000000 ;
			15'h0000629D : data <= 8'b00000000 ;
			15'h0000629E : data <= 8'b00000000 ;
			15'h0000629F : data <= 8'b00000000 ;
			15'h000062A0 : data <= 8'b00000000 ;
			15'h000062A1 : data <= 8'b00000000 ;
			15'h000062A2 : data <= 8'b00000000 ;
			15'h000062A3 : data <= 8'b00000000 ;
			15'h000062A4 : data <= 8'b00000000 ;
			15'h000062A5 : data <= 8'b00000000 ;
			15'h000062A6 : data <= 8'b00000000 ;
			15'h000062A7 : data <= 8'b00000000 ;
			15'h000062A8 : data <= 8'b00000000 ;
			15'h000062A9 : data <= 8'b00000000 ;
			15'h000062AA : data <= 8'b00000000 ;
			15'h000062AB : data <= 8'b00000000 ;
			15'h000062AC : data <= 8'b00000000 ;
			15'h000062AD : data <= 8'b00000000 ;
			15'h000062AE : data <= 8'b00000000 ;
			15'h000062AF : data <= 8'b00000000 ;
			15'h000062B0 : data <= 8'b00000000 ;
			15'h000062B1 : data <= 8'b00000000 ;
			15'h000062B2 : data <= 8'b00000000 ;
			15'h000062B3 : data <= 8'b00000000 ;
			15'h000062B4 : data <= 8'b00000000 ;
			15'h000062B5 : data <= 8'b00000000 ;
			15'h000062B6 : data <= 8'b00000000 ;
			15'h000062B7 : data <= 8'b00000000 ;
			15'h000062B8 : data <= 8'b00000000 ;
			15'h000062B9 : data <= 8'b00000000 ;
			15'h000062BA : data <= 8'b00000000 ;
			15'h000062BB : data <= 8'b00000000 ;
			15'h000062BC : data <= 8'b00000000 ;
			15'h000062BD : data <= 8'b00000000 ;
			15'h000062BE : data <= 8'b00000000 ;
			15'h000062BF : data <= 8'b00000000 ;
			15'h000062C0 : data <= 8'b00000000 ;
			15'h000062C1 : data <= 8'b00000000 ;
			15'h000062C2 : data <= 8'b00000000 ;
			15'h000062C3 : data <= 8'b00000000 ;
			15'h000062C4 : data <= 8'b00000000 ;
			15'h000062C5 : data <= 8'b00000000 ;
			15'h000062C6 : data <= 8'b00000000 ;
			15'h000062C7 : data <= 8'b00000000 ;
			15'h000062C8 : data <= 8'b00000000 ;
			15'h000062C9 : data <= 8'b00000000 ;
			15'h000062CA : data <= 8'b00000000 ;
			15'h000062CB : data <= 8'b00000000 ;
			15'h000062CC : data <= 8'b00000000 ;
			15'h000062CD : data <= 8'b00000000 ;
			15'h000062CE : data <= 8'b00000000 ;
			15'h000062CF : data <= 8'b00000000 ;
			15'h000062D0 : data <= 8'b00000000 ;
			15'h000062D1 : data <= 8'b00000000 ;
			15'h000062D2 : data <= 8'b00000000 ;
			15'h000062D3 : data <= 8'b00000000 ;
			15'h000062D4 : data <= 8'b00000000 ;
			15'h000062D5 : data <= 8'b00000000 ;
			15'h000062D6 : data <= 8'b00000000 ;
			15'h000062D7 : data <= 8'b00000000 ;
			15'h000062D8 : data <= 8'b00000000 ;
			15'h000062D9 : data <= 8'b00000000 ;
			15'h000062DA : data <= 8'b00000000 ;
			15'h000062DB : data <= 8'b00000000 ;
			15'h000062DC : data <= 8'b00000000 ;
			15'h000062DD : data <= 8'b00000000 ;
			15'h000062DE : data <= 8'b00000000 ;
			15'h000062DF : data <= 8'b00000000 ;
			15'h000062E0 : data <= 8'b00000000 ;
			15'h000062E1 : data <= 8'b00000000 ;
			15'h000062E2 : data <= 8'b00000000 ;
			15'h000062E3 : data <= 8'b00000000 ;
			15'h000062E4 : data <= 8'b00000000 ;
			15'h000062E5 : data <= 8'b00000000 ;
			15'h000062E6 : data <= 8'b00000000 ;
			15'h000062E7 : data <= 8'b00000000 ;
			15'h000062E8 : data <= 8'b00000000 ;
			15'h000062E9 : data <= 8'b00000000 ;
			15'h000062EA : data <= 8'b00000000 ;
			15'h000062EB : data <= 8'b00000000 ;
			15'h000062EC : data <= 8'b00000000 ;
			15'h000062ED : data <= 8'b00000000 ;
			15'h000062EE : data <= 8'b00000000 ;
			15'h000062EF : data <= 8'b00000000 ;
			15'h000062F0 : data <= 8'b00000000 ;
			15'h000062F1 : data <= 8'b00000000 ;
			15'h000062F2 : data <= 8'b00000000 ;
			15'h000062F3 : data <= 8'b00000000 ;
			15'h000062F4 : data <= 8'b00000000 ;
			15'h000062F5 : data <= 8'b00000000 ;
			15'h000062F6 : data <= 8'b00000000 ;
			15'h000062F7 : data <= 8'b00000000 ;
			15'h000062F8 : data <= 8'b00000000 ;
			15'h000062F9 : data <= 8'b00000000 ;
			15'h000062FA : data <= 8'b00000000 ;
			15'h000062FB : data <= 8'b00000000 ;
			15'h000062FC : data <= 8'b00000000 ;
			15'h000062FD : data <= 8'b00000000 ;
			15'h000062FE : data <= 8'b00000000 ;
			15'h000062FF : data <= 8'b00000000 ;
			15'h00006300 : data <= 8'b00000000 ;
			15'h00006301 : data <= 8'b00000000 ;
			15'h00006302 : data <= 8'b00000000 ;
			15'h00006303 : data <= 8'b00000000 ;
			15'h00006304 : data <= 8'b00000000 ;
			15'h00006305 : data <= 8'b00000000 ;
			15'h00006306 : data <= 8'b00000000 ;
			15'h00006307 : data <= 8'b00000000 ;
			15'h00006308 : data <= 8'b00000000 ;
			15'h00006309 : data <= 8'b00000000 ;
			15'h0000630A : data <= 8'b00000000 ;
			15'h0000630B : data <= 8'b00000000 ;
			15'h0000630C : data <= 8'b00000000 ;
			15'h0000630D : data <= 8'b00000000 ;
			15'h0000630E : data <= 8'b00000000 ;
			15'h0000630F : data <= 8'b00000000 ;
			15'h00006310 : data <= 8'b00000000 ;
			15'h00006311 : data <= 8'b00000000 ;
			15'h00006312 : data <= 8'b00000000 ;
			15'h00006313 : data <= 8'b00000000 ;
			15'h00006314 : data <= 8'b00000000 ;
			15'h00006315 : data <= 8'b00000000 ;
			15'h00006316 : data <= 8'b00000000 ;
			15'h00006317 : data <= 8'b00000000 ;
			15'h00006318 : data <= 8'b00000000 ;
			15'h00006319 : data <= 8'b00000000 ;
			15'h0000631A : data <= 8'b00000000 ;
			15'h0000631B : data <= 8'b00000000 ;
			15'h0000631C : data <= 8'b00000000 ;
			15'h0000631D : data <= 8'b00000000 ;
			15'h0000631E : data <= 8'b00000000 ;
			15'h0000631F : data <= 8'b00000000 ;
			15'h00006320 : data <= 8'b00000000 ;
			15'h00006321 : data <= 8'b00000000 ;
			15'h00006322 : data <= 8'b00000000 ;
			15'h00006323 : data <= 8'b00000000 ;
			15'h00006324 : data <= 8'b00000000 ;
			15'h00006325 : data <= 8'b00000000 ;
			15'h00006326 : data <= 8'b00000000 ;
			15'h00006327 : data <= 8'b00000000 ;
			15'h00006328 : data <= 8'b00000000 ;
			15'h00006329 : data <= 8'b00000000 ;
			15'h0000632A : data <= 8'b00000000 ;
			15'h0000632B : data <= 8'b00000000 ;
			15'h0000632C : data <= 8'b00000000 ;
			15'h0000632D : data <= 8'b00000000 ;
			15'h0000632E : data <= 8'b00000000 ;
			15'h0000632F : data <= 8'b00000000 ;
			15'h00006330 : data <= 8'b00000000 ;
			15'h00006331 : data <= 8'b00000000 ;
			15'h00006332 : data <= 8'b00000000 ;
			15'h00006333 : data <= 8'b00000000 ;
			15'h00006334 : data <= 8'b00000000 ;
			15'h00006335 : data <= 8'b00000000 ;
			15'h00006336 : data <= 8'b00000000 ;
			15'h00006337 : data <= 8'b00000000 ;
			15'h00006338 : data <= 8'b00000000 ;
			15'h00006339 : data <= 8'b00000000 ;
			15'h0000633A : data <= 8'b00000000 ;
			15'h0000633B : data <= 8'b00000000 ;
			15'h0000633C : data <= 8'b00000000 ;
			15'h0000633D : data <= 8'b00000000 ;
			15'h0000633E : data <= 8'b00000000 ;
			15'h0000633F : data <= 8'b00000000 ;
			15'h00006340 : data <= 8'b00000000 ;
			15'h00006341 : data <= 8'b00000000 ;
			15'h00006342 : data <= 8'b00000000 ;
			15'h00006343 : data <= 8'b00000000 ;
			15'h00006344 : data <= 8'b00000000 ;
			15'h00006345 : data <= 8'b00000000 ;
			15'h00006346 : data <= 8'b00000000 ;
			15'h00006347 : data <= 8'b00000000 ;
			15'h00006348 : data <= 8'b00000000 ;
			15'h00006349 : data <= 8'b00000000 ;
			15'h0000634A : data <= 8'b00000000 ;
			15'h0000634B : data <= 8'b00000000 ;
			15'h0000634C : data <= 8'b00000000 ;
			15'h0000634D : data <= 8'b00000000 ;
			15'h0000634E : data <= 8'b00000000 ;
			15'h0000634F : data <= 8'b00000000 ;
			15'h00006350 : data <= 8'b00000000 ;
			15'h00006351 : data <= 8'b00000000 ;
			15'h00006352 : data <= 8'b00000000 ;
			15'h00006353 : data <= 8'b00000000 ;
			15'h00006354 : data <= 8'b00000000 ;
			15'h00006355 : data <= 8'b00000000 ;
			15'h00006356 : data <= 8'b00000000 ;
			15'h00006357 : data <= 8'b00000000 ;
			15'h00006358 : data <= 8'b00000000 ;
			15'h00006359 : data <= 8'b00000000 ;
			15'h0000635A : data <= 8'b00000000 ;
			15'h0000635B : data <= 8'b00000000 ;
			15'h0000635C : data <= 8'b00000000 ;
			15'h0000635D : data <= 8'b00000000 ;
			15'h0000635E : data <= 8'b00000000 ;
			15'h0000635F : data <= 8'b00000000 ;
			15'h00006360 : data <= 8'b00000000 ;
			15'h00006361 : data <= 8'b00000000 ;
			15'h00006362 : data <= 8'b00000000 ;
			15'h00006363 : data <= 8'b00000000 ;
			15'h00006364 : data <= 8'b00000000 ;
			15'h00006365 : data <= 8'b00000000 ;
			15'h00006366 : data <= 8'b00000000 ;
			15'h00006367 : data <= 8'b00000000 ;
			15'h00006368 : data <= 8'b00000000 ;
			15'h00006369 : data <= 8'b00000000 ;
			15'h0000636A : data <= 8'b00000000 ;
			15'h0000636B : data <= 8'b00000000 ;
			15'h0000636C : data <= 8'b00000000 ;
			15'h0000636D : data <= 8'b00000000 ;
			15'h0000636E : data <= 8'b00000000 ;
			15'h0000636F : data <= 8'b00000000 ;
			15'h00006370 : data <= 8'b00000000 ;
			15'h00006371 : data <= 8'b00000000 ;
			15'h00006372 : data <= 8'b00000000 ;
			15'h00006373 : data <= 8'b00000000 ;
			15'h00006374 : data <= 8'b00000000 ;
			15'h00006375 : data <= 8'b00000000 ;
			15'h00006376 : data <= 8'b00000000 ;
			15'h00006377 : data <= 8'b00000000 ;
			15'h00006378 : data <= 8'b00000000 ;
			15'h00006379 : data <= 8'b00000000 ;
			15'h0000637A : data <= 8'b00000000 ;
			15'h0000637B : data <= 8'b00000000 ;
			15'h0000637C : data <= 8'b00000000 ;
			15'h0000637D : data <= 8'b00000000 ;
			15'h0000637E : data <= 8'b00000000 ;
			15'h0000637F : data <= 8'b00000000 ;
			15'h00006380 : data <= 8'b00000000 ;
			15'h00006381 : data <= 8'b00000000 ;
			15'h00006382 : data <= 8'b00000000 ;
			15'h00006383 : data <= 8'b00000000 ;
			15'h00006384 : data <= 8'b00000000 ;
			15'h00006385 : data <= 8'b00000000 ;
			15'h00006386 : data <= 8'b00000000 ;
			15'h00006387 : data <= 8'b00000000 ;
			15'h00006388 : data <= 8'b00000000 ;
			15'h00006389 : data <= 8'b00000000 ;
			15'h0000638A : data <= 8'b00000000 ;
			15'h0000638B : data <= 8'b00000000 ;
			15'h0000638C : data <= 8'b00000000 ;
			15'h0000638D : data <= 8'b00000000 ;
			15'h0000638E : data <= 8'b00000000 ;
			15'h0000638F : data <= 8'b00000000 ;
			15'h00006390 : data <= 8'b00000000 ;
			15'h00006391 : data <= 8'b00000000 ;
			15'h00006392 : data <= 8'b00000000 ;
			15'h00006393 : data <= 8'b00000000 ;
			15'h00006394 : data <= 8'b00000000 ;
			15'h00006395 : data <= 8'b00000000 ;
			15'h00006396 : data <= 8'b00000000 ;
			15'h00006397 : data <= 8'b00000000 ;
			15'h00006398 : data <= 8'b00000000 ;
			15'h00006399 : data <= 8'b00000000 ;
			15'h0000639A : data <= 8'b00000000 ;
			15'h0000639B : data <= 8'b00000000 ;
			15'h0000639C : data <= 8'b00000000 ;
			15'h0000639D : data <= 8'b00000000 ;
			15'h0000639E : data <= 8'b00000000 ;
			15'h0000639F : data <= 8'b00000000 ;
			15'h000063A0 : data <= 8'b00000000 ;
			15'h000063A1 : data <= 8'b00000000 ;
			15'h000063A2 : data <= 8'b00000000 ;
			15'h000063A3 : data <= 8'b00000000 ;
			15'h000063A4 : data <= 8'b00000000 ;
			15'h000063A5 : data <= 8'b00000000 ;
			15'h000063A6 : data <= 8'b00000000 ;
			15'h000063A7 : data <= 8'b00000000 ;
			15'h000063A8 : data <= 8'b00000000 ;
			15'h000063A9 : data <= 8'b00000000 ;
			15'h000063AA : data <= 8'b00000000 ;
			15'h000063AB : data <= 8'b00000000 ;
			15'h000063AC : data <= 8'b00000000 ;
			15'h000063AD : data <= 8'b00000000 ;
			15'h000063AE : data <= 8'b00000000 ;
			15'h000063AF : data <= 8'b00000000 ;
			15'h000063B0 : data <= 8'b00000000 ;
			15'h000063B1 : data <= 8'b00000000 ;
			15'h000063B2 : data <= 8'b00000000 ;
			15'h000063B3 : data <= 8'b00000000 ;
			15'h000063B4 : data <= 8'b00000000 ;
			15'h000063B5 : data <= 8'b00000000 ;
			15'h000063B6 : data <= 8'b00000000 ;
			15'h000063B7 : data <= 8'b00000000 ;
			15'h000063B8 : data <= 8'b00000000 ;
			15'h000063B9 : data <= 8'b00000000 ;
			15'h000063BA : data <= 8'b00000000 ;
			15'h000063BB : data <= 8'b00000000 ;
			15'h000063BC : data <= 8'b00000000 ;
			15'h000063BD : data <= 8'b00000000 ;
			15'h000063BE : data <= 8'b00000000 ;
			15'h000063BF : data <= 8'b00000000 ;
			15'h000063C0 : data <= 8'b00000000 ;
			15'h000063C1 : data <= 8'b00000000 ;
			15'h000063C2 : data <= 8'b00000000 ;
			15'h000063C3 : data <= 8'b00000000 ;
			15'h000063C4 : data <= 8'b00000000 ;
			15'h000063C5 : data <= 8'b00000000 ;
			15'h000063C6 : data <= 8'b00000000 ;
			15'h000063C7 : data <= 8'b00000000 ;
			15'h000063C8 : data <= 8'b00000000 ;
			15'h000063C9 : data <= 8'b00000000 ;
			15'h000063CA : data <= 8'b00000000 ;
			15'h000063CB : data <= 8'b00000000 ;
			15'h000063CC : data <= 8'b00000000 ;
			15'h000063CD : data <= 8'b00000000 ;
			15'h000063CE : data <= 8'b00000000 ;
			15'h000063CF : data <= 8'b00000000 ;
			15'h000063D0 : data <= 8'b00000000 ;
			15'h000063D1 : data <= 8'b00000000 ;
			15'h000063D2 : data <= 8'b00000000 ;
			15'h000063D3 : data <= 8'b00000000 ;
			15'h000063D4 : data <= 8'b00000000 ;
			15'h000063D5 : data <= 8'b00000000 ;
			15'h000063D6 : data <= 8'b00000000 ;
			15'h000063D7 : data <= 8'b00000000 ;
			15'h000063D8 : data <= 8'b00000000 ;
			15'h000063D9 : data <= 8'b00000000 ;
			15'h000063DA : data <= 8'b00000000 ;
			15'h000063DB : data <= 8'b00000000 ;
			15'h000063DC : data <= 8'b00000000 ;
			15'h000063DD : data <= 8'b00000000 ;
			15'h000063DE : data <= 8'b00000000 ;
			15'h000063DF : data <= 8'b00000000 ;
			15'h000063E0 : data <= 8'b00000000 ;
			15'h000063E1 : data <= 8'b00000000 ;
			15'h000063E2 : data <= 8'b00000000 ;
			15'h000063E3 : data <= 8'b00000000 ;
			15'h000063E4 : data <= 8'b00000000 ;
			15'h000063E5 : data <= 8'b00000000 ;
			15'h000063E6 : data <= 8'b00000000 ;
			15'h000063E7 : data <= 8'b00000000 ;
			15'h000063E8 : data <= 8'b00000000 ;
			15'h000063E9 : data <= 8'b00000000 ;
			15'h000063EA : data <= 8'b00000000 ;
			15'h000063EB : data <= 8'b00000000 ;
			15'h000063EC : data <= 8'b00000000 ;
			15'h000063ED : data <= 8'b00000000 ;
			15'h000063EE : data <= 8'b00000000 ;
			15'h000063EF : data <= 8'b00000000 ;
			15'h000063F0 : data <= 8'b00000000 ;
			15'h000063F1 : data <= 8'b00000000 ;
			15'h000063F2 : data <= 8'b00000000 ;
			15'h000063F3 : data <= 8'b00000000 ;
			15'h000063F4 : data <= 8'b00000000 ;
			15'h000063F5 : data <= 8'b00000000 ;
			15'h000063F6 : data <= 8'b00000000 ;
			15'h000063F7 : data <= 8'b00000000 ;
			15'h000063F8 : data <= 8'b00000000 ;
			15'h000063F9 : data <= 8'b00000000 ;
			15'h000063FA : data <= 8'b00000000 ;
			15'h000063FB : data <= 8'b00000000 ;
			15'h000063FC : data <= 8'b00000000 ;
			15'h000063FD : data <= 8'b00000000 ;
			15'h000063FE : data <= 8'b00000000 ;
			15'h000063FF : data <= 8'b00000000 ;
			15'h00006400 : data <= 8'b00000000 ;
			15'h00006401 : data <= 8'b00000000 ;
			15'h00006402 : data <= 8'b00000000 ;
			15'h00006403 : data <= 8'b00000000 ;
			15'h00006404 : data <= 8'b00000000 ;
			15'h00006405 : data <= 8'b00000000 ;
			15'h00006406 : data <= 8'b00000000 ;
			15'h00006407 : data <= 8'b00000000 ;
			15'h00006408 : data <= 8'b00000000 ;
			15'h00006409 : data <= 8'b00000000 ;
			15'h0000640A : data <= 8'b00000000 ;
			15'h0000640B : data <= 8'b00000000 ;
			15'h0000640C : data <= 8'b00000000 ;
			15'h0000640D : data <= 8'b00000000 ;
			15'h0000640E : data <= 8'b00000000 ;
			15'h0000640F : data <= 8'b00000000 ;
			15'h00006410 : data <= 8'b00000000 ;
			15'h00006411 : data <= 8'b00000000 ;
			15'h00006412 : data <= 8'b00000000 ;
			15'h00006413 : data <= 8'b00000000 ;
			15'h00006414 : data <= 8'b00000000 ;
			15'h00006415 : data <= 8'b00000000 ;
			15'h00006416 : data <= 8'b00000000 ;
			15'h00006417 : data <= 8'b00000000 ;
			15'h00006418 : data <= 8'b00000000 ;
			15'h00006419 : data <= 8'b00000000 ;
			15'h0000641A : data <= 8'b00000000 ;
			15'h0000641B : data <= 8'b00000000 ;
			15'h0000641C : data <= 8'b00000000 ;
			15'h0000641D : data <= 8'b00000000 ;
			15'h0000641E : data <= 8'b00000000 ;
			15'h0000641F : data <= 8'b00000000 ;
			15'h00006420 : data <= 8'b00000000 ;
			15'h00006421 : data <= 8'b00000000 ;
			15'h00006422 : data <= 8'b00000000 ;
			15'h00006423 : data <= 8'b00000000 ;
			15'h00006424 : data <= 8'b00000000 ;
			15'h00006425 : data <= 8'b00000000 ;
			15'h00006426 : data <= 8'b00000000 ;
			15'h00006427 : data <= 8'b00000000 ;
			15'h00006428 : data <= 8'b00000000 ;
			15'h00006429 : data <= 8'b00000000 ;
			15'h0000642A : data <= 8'b00000000 ;
			15'h0000642B : data <= 8'b00000000 ;
			15'h0000642C : data <= 8'b00000000 ;
			15'h0000642D : data <= 8'b00000000 ;
			15'h0000642E : data <= 8'b00000000 ;
			15'h0000642F : data <= 8'b00000000 ;
			15'h00006430 : data <= 8'b00000000 ;
			15'h00006431 : data <= 8'b00000000 ;
			15'h00006432 : data <= 8'b00000000 ;
			15'h00006433 : data <= 8'b00000000 ;
			15'h00006434 : data <= 8'b00000000 ;
			15'h00006435 : data <= 8'b00000000 ;
			15'h00006436 : data <= 8'b00000000 ;
			15'h00006437 : data <= 8'b00000000 ;
			15'h00006438 : data <= 8'b00000000 ;
			15'h00006439 : data <= 8'b00000000 ;
			15'h0000643A : data <= 8'b00000000 ;
			15'h0000643B : data <= 8'b00000000 ;
			15'h0000643C : data <= 8'b00000000 ;
			15'h0000643D : data <= 8'b00000000 ;
			15'h0000643E : data <= 8'b00000000 ;
			15'h0000643F : data <= 8'b00000000 ;
			15'h00006440 : data <= 8'b00000000 ;
			15'h00006441 : data <= 8'b00000000 ;
			15'h00006442 : data <= 8'b00000000 ;
			15'h00006443 : data <= 8'b00000000 ;
			15'h00006444 : data <= 8'b00000000 ;
			15'h00006445 : data <= 8'b00000000 ;
			15'h00006446 : data <= 8'b00000000 ;
			15'h00006447 : data <= 8'b00000000 ;
			15'h00006448 : data <= 8'b00000000 ;
			15'h00006449 : data <= 8'b00000000 ;
			15'h0000644A : data <= 8'b00000000 ;
			15'h0000644B : data <= 8'b00000000 ;
			15'h0000644C : data <= 8'b00000000 ;
			15'h0000644D : data <= 8'b00000000 ;
			15'h0000644E : data <= 8'b00000000 ;
			15'h0000644F : data <= 8'b00000000 ;
			15'h00006450 : data <= 8'b00000000 ;
			15'h00006451 : data <= 8'b00000000 ;
			15'h00006452 : data <= 8'b00000000 ;
			15'h00006453 : data <= 8'b00000000 ;
			15'h00006454 : data <= 8'b00000000 ;
			15'h00006455 : data <= 8'b00000000 ;
			15'h00006456 : data <= 8'b00000000 ;
			15'h00006457 : data <= 8'b00000000 ;
			15'h00006458 : data <= 8'b00000000 ;
			15'h00006459 : data <= 8'b00000000 ;
			15'h0000645A : data <= 8'b00000000 ;
			15'h0000645B : data <= 8'b00000000 ;
			15'h0000645C : data <= 8'b00000000 ;
			15'h0000645D : data <= 8'b00000000 ;
			15'h0000645E : data <= 8'b00000000 ;
			15'h0000645F : data <= 8'b00000000 ;
			15'h00006460 : data <= 8'b00000000 ;
			15'h00006461 : data <= 8'b00000000 ;
			15'h00006462 : data <= 8'b00000000 ;
			15'h00006463 : data <= 8'b00000000 ;
			15'h00006464 : data <= 8'b00000000 ;
			15'h00006465 : data <= 8'b00000000 ;
			15'h00006466 : data <= 8'b00000000 ;
			15'h00006467 : data <= 8'b00000000 ;
			15'h00006468 : data <= 8'b00000000 ;
			15'h00006469 : data <= 8'b00000000 ;
			15'h0000646A : data <= 8'b00000000 ;
			15'h0000646B : data <= 8'b00000000 ;
			15'h0000646C : data <= 8'b00000000 ;
			15'h0000646D : data <= 8'b00000000 ;
			15'h0000646E : data <= 8'b00000000 ;
			15'h0000646F : data <= 8'b00000000 ;
			15'h00006470 : data <= 8'b00000000 ;
			15'h00006471 : data <= 8'b00000000 ;
			15'h00006472 : data <= 8'b00000000 ;
			15'h00006473 : data <= 8'b00000000 ;
			15'h00006474 : data <= 8'b00000000 ;
			15'h00006475 : data <= 8'b00000000 ;
			15'h00006476 : data <= 8'b00000000 ;
			15'h00006477 : data <= 8'b00000000 ;
			15'h00006478 : data <= 8'b00000000 ;
			15'h00006479 : data <= 8'b00000000 ;
			15'h0000647A : data <= 8'b00000000 ;
			15'h0000647B : data <= 8'b00000000 ;
			15'h0000647C : data <= 8'b00000000 ;
			15'h0000647D : data <= 8'b00000000 ;
			15'h0000647E : data <= 8'b00000000 ;
			15'h0000647F : data <= 8'b00000000 ;
			15'h00006480 : data <= 8'b00000000 ;
			15'h00006481 : data <= 8'b00000000 ;
			15'h00006482 : data <= 8'b00000000 ;
			15'h00006483 : data <= 8'b00000000 ;
			15'h00006484 : data <= 8'b00000000 ;
			15'h00006485 : data <= 8'b00000000 ;
			15'h00006486 : data <= 8'b00000000 ;
			15'h00006487 : data <= 8'b00000000 ;
			15'h00006488 : data <= 8'b00000000 ;
			15'h00006489 : data <= 8'b00000000 ;
			15'h0000648A : data <= 8'b00000000 ;
			15'h0000648B : data <= 8'b00000000 ;
			15'h0000648C : data <= 8'b00000000 ;
			15'h0000648D : data <= 8'b00000000 ;
			15'h0000648E : data <= 8'b00000000 ;
			15'h0000648F : data <= 8'b00000000 ;
			15'h00006490 : data <= 8'b00000000 ;
			15'h00006491 : data <= 8'b00000000 ;
			15'h00006492 : data <= 8'b00000000 ;
			15'h00006493 : data <= 8'b00000000 ;
			15'h00006494 : data <= 8'b00000000 ;
			15'h00006495 : data <= 8'b00000000 ;
			15'h00006496 : data <= 8'b00000000 ;
			15'h00006497 : data <= 8'b00000000 ;
			15'h00006498 : data <= 8'b00000000 ;
			15'h00006499 : data <= 8'b00000000 ;
			15'h0000649A : data <= 8'b00000000 ;
			15'h0000649B : data <= 8'b00000000 ;
			15'h0000649C : data <= 8'b00000000 ;
			15'h0000649D : data <= 8'b00000000 ;
			15'h0000649E : data <= 8'b00000000 ;
			15'h0000649F : data <= 8'b00000000 ;
			15'h000064A0 : data <= 8'b00000000 ;
			15'h000064A1 : data <= 8'b00000000 ;
			15'h000064A2 : data <= 8'b00000000 ;
			15'h000064A3 : data <= 8'b00000000 ;
			15'h000064A4 : data <= 8'b00000000 ;
			15'h000064A5 : data <= 8'b00000000 ;
			15'h000064A6 : data <= 8'b00000000 ;
			15'h000064A7 : data <= 8'b00000000 ;
			15'h000064A8 : data <= 8'b00000000 ;
			15'h000064A9 : data <= 8'b00000000 ;
			15'h000064AA : data <= 8'b00000000 ;
			15'h000064AB : data <= 8'b00000000 ;
			15'h000064AC : data <= 8'b00000000 ;
			15'h000064AD : data <= 8'b00000000 ;
			15'h000064AE : data <= 8'b00000000 ;
			15'h000064AF : data <= 8'b00000000 ;
			15'h000064B0 : data <= 8'b00000000 ;
			15'h000064B1 : data <= 8'b00000000 ;
			15'h000064B2 : data <= 8'b00000000 ;
			15'h000064B3 : data <= 8'b00000000 ;
			15'h000064B4 : data <= 8'b00000000 ;
			15'h000064B5 : data <= 8'b00000000 ;
			15'h000064B6 : data <= 8'b00000000 ;
			15'h000064B7 : data <= 8'b00000000 ;
			15'h000064B8 : data <= 8'b00000000 ;
			15'h000064B9 : data <= 8'b00000000 ;
			15'h000064BA : data <= 8'b00000000 ;
			15'h000064BB : data <= 8'b00000000 ;
			15'h000064BC : data <= 8'b00000000 ;
			15'h000064BD : data <= 8'b00000000 ;
			15'h000064BE : data <= 8'b00000000 ;
			15'h000064BF : data <= 8'b00000000 ;
			15'h000064C0 : data <= 8'b00000000 ;
			15'h000064C1 : data <= 8'b00000000 ;
			15'h000064C2 : data <= 8'b00000000 ;
			15'h000064C3 : data <= 8'b00000000 ;
			15'h000064C4 : data <= 8'b00000000 ;
			15'h000064C5 : data <= 8'b00000000 ;
			15'h000064C6 : data <= 8'b00000000 ;
			15'h000064C7 : data <= 8'b00000000 ;
			15'h000064C8 : data <= 8'b00000000 ;
			15'h000064C9 : data <= 8'b00000000 ;
			15'h000064CA : data <= 8'b00000000 ;
			15'h000064CB : data <= 8'b00000000 ;
			15'h000064CC : data <= 8'b00000000 ;
			15'h000064CD : data <= 8'b00000000 ;
			15'h000064CE : data <= 8'b00000000 ;
			15'h000064CF : data <= 8'b00000000 ;
			15'h000064D0 : data <= 8'b00000000 ;
			15'h000064D1 : data <= 8'b00000000 ;
			15'h000064D2 : data <= 8'b00000000 ;
			15'h000064D3 : data <= 8'b00000000 ;
			15'h000064D4 : data <= 8'b00000000 ;
			15'h000064D5 : data <= 8'b00000000 ;
			15'h000064D6 : data <= 8'b00000000 ;
			15'h000064D7 : data <= 8'b00000000 ;
			15'h000064D8 : data <= 8'b00000000 ;
			15'h000064D9 : data <= 8'b00000000 ;
			15'h000064DA : data <= 8'b00000000 ;
			15'h000064DB : data <= 8'b00000000 ;
			15'h000064DC : data <= 8'b00000000 ;
			15'h000064DD : data <= 8'b00000000 ;
			15'h000064DE : data <= 8'b00000000 ;
			15'h000064DF : data <= 8'b00000000 ;
			15'h000064E0 : data <= 8'b00000000 ;
			15'h000064E1 : data <= 8'b00000000 ;
			15'h000064E2 : data <= 8'b00000000 ;
			15'h000064E3 : data <= 8'b00000000 ;
			15'h000064E4 : data <= 8'b00000000 ;
			15'h000064E5 : data <= 8'b00000000 ;
			15'h000064E6 : data <= 8'b00000000 ;
			15'h000064E7 : data <= 8'b00000000 ;
			15'h000064E8 : data <= 8'b00000000 ;
			15'h000064E9 : data <= 8'b00000000 ;
			15'h000064EA : data <= 8'b00000000 ;
			15'h000064EB : data <= 8'b00000000 ;
			15'h000064EC : data <= 8'b00000000 ;
			15'h000064ED : data <= 8'b00000000 ;
			15'h000064EE : data <= 8'b00000000 ;
			15'h000064EF : data <= 8'b00000000 ;
			15'h000064F0 : data <= 8'b00000000 ;
			15'h000064F1 : data <= 8'b00000000 ;
			15'h000064F2 : data <= 8'b00000000 ;
			15'h000064F3 : data <= 8'b00000000 ;
			15'h000064F4 : data <= 8'b00000000 ;
			15'h000064F5 : data <= 8'b00000000 ;
			15'h000064F6 : data <= 8'b00000000 ;
			15'h000064F7 : data <= 8'b00000000 ;
			15'h000064F8 : data <= 8'b00000000 ;
			15'h000064F9 : data <= 8'b00000000 ;
			15'h000064FA : data <= 8'b00000000 ;
			15'h000064FB : data <= 8'b00000000 ;
			15'h000064FC : data <= 8'b00000000 ;
			15'h000064FD : data <= 8'b00000000 ;
			15'h000064FE : data <= 8'b00000000 ;
			15'h000064FF : data <= 8'b00000000 ;
			15'h00006500 : data <= 8'b00000000 ;
			15'h00006501 : data <= 8'b00000000 ;
			15'h00006502 : data <= 8'b00000000 ;
			15'h00006503 : data <= 8'b00000000 ;
			15'h00006504 : data <= 8'b00000000 ;
			15'h00006505 : data <= 8'b00000000 ;
			15'h00006506 : data <= 8'b00000000 ;
			15'h00006507 : data <= 8'b00000000 ;
			15'h00006508 : data <= 8'b00000000 ;
			15'h00006509 : data <= 8'b00000000 ;
			15'h0000650A : data <= 8'b00000000 ;
			15'h0000650B : data <= 8'b00000000 ;
			15'h0000650C : data <= 8'b00000000 ;
			15'h0000650D : data <= 8'b00000000 ;
			15'h0000650E : data <= 8'b00000000 ;
			15'h0000650F : data <= 8'b00000000 ;
			15'h00006510 : data <= 8'b00000000 ;
			15'h00006511 : data <= 8'b00000000 ;
			15'h00006512 : data <= 8'b00000000 ;
			15'h00006513 : data <= 8'b00000000 ;
			15'h00006514 : data <= 8'b00000000 ;
			15'h00006515 : data <= 8'b00000000 ;
			15'h00006516 : data <= 8'b00000000 ;
			15'h00006517 : data <= 8'b00000000 ;
			15'h00006518 : data <= 8'b00000000 ;
			15'h00006519 : data <= 8'b00000000 ;
			15'h0000651A : data <= 8'b00000000 ;
			15'h0000651B : data <= 8'b00000000 ;
			15'h0000651C : data <= 8'b00000000 ;
			15'h0000651D : data <= 8'b00000000 ;
			15'h0000651E : data <= 8'b00000000 ;
			15'h0000651F : data <= 8'b00000000 ;
			15'h00006520 : data <= 8'b00000000 ;
			15'h00006521 : data <= 8'b00000000 ;
			15'h00006522 : data <= 8'b00000000 ;
			15'h00006523 : data <= 8'b00000000 ;
			15'h00006524 : data <= 8'b00000000 ;
			15'h00006525 : data <= 8'b00000000 ;
			15'h00006526 : data <= 8'b00000000 ;
			15'h00006527 : data <= 8'b00000000 ;
			15'h00006528 : data <= 8'b00000000 ;
			15'h00006529 : data <= 8'b00000000 ;
			15'h0000652A : data <= 8'b00000000 ;
			15'h0000652B : data <= 8'b00000000 ;
			15'h0000652C : data <= 8'b00000000 ;
			15'h0000652D : data <= 8'b00000000 ;
			15'h0000652E : data <= 8'b00000000 ;
			15'h0000652F : data <= 8'b00000000 ;
			15'h00006530 : data <= 8'b00000000 ;
			15'h00006531 : data <= 8'b00000000 ;
			15'h00006532 : data <= 8'b00000000 ;
			15'h00006533 : data <= 8'b00000000 ;
			15'h00006534 : data <= 8'b00000000 ;
			15'h00006535 : data <= 8'b00000000 ;
			15'h00006536 : data <= 8'b00000000 ;
			15'h00006537 : data <= 8'b00000000 ;
			15'h00006538 : data <= 8'b00000000 ;
			15'h00006539 : data <= 8'b00000000 ;
			15'h0000653A : data <= 8'b00000000 ;
			15'h0000653B : data <= 8'b00000000 ;
			15'h0000653C : data <= 8'b00000000 ;
			15'h0000653D : data <= 8'b00000000 ;
			15'h0000653E : data <= 8'b00000000 ;
			15'h0000653F : data <= 8'b00000000 ;
			15'h00006540 : data <= 8'b00000000 ;
			15'h00006541 : data <= 8'b00000000 ;
			15'h00006542 : data <= 8'b00000000 ;
			15'h00006543 : data <= 8'b00000000 ;
			15'h00006544 : data <= 8'b00000000 ;
			15'h00006545 : data <= 8'b00000000 ;
			15'h00006546 : data <= 8'b00000000 ;
			15'h00006547 : data <= 8'b00000000 ;
			15'h00006548 : data <= 8'b00000000 ;
			15'h00006549 : data <= 8'b00000000 ;
			15'h0000654A : data <= 8'b00000000 ;
			15'h0000654B : data <= 8'b00000000 ;
			15'h0000654C : data <= 8'b00000000 ;
			15'h0000654D : data <= 8'b00000000 ;
			15'h0000654E : data <= 8'b00000000 ;
			15'h0000654F : data <= 8'b00000000 ;
			15'h00006550 : data <= 8'b00000000 ;
			15'h00006551 : data <= 8'b00000000 ;
			15'h00006552 : data <= 8'b00000000 ;
			15'h00006553 : data <= 8'b00000000 ;
			15'h00006554 : data <= 8'b00000000 ;
			15'h00006555 : data <= 8'b00000000 ;
			15'h00006556 : data <= 8'b00000000 ;
			15'h00006557 : data <= 8'b00000000 ;
			15'h00006558 : data <= 8'b00000000 ;
			15'h00006559 : data <= 8'b00000000 ;
			15'h0000655A : data <= 8'b00000000 ;
			15'h0000655B : data <= 8'b00000000 ;
			15'h0000655C : data <= 8'b00000000 ;
			15'h0000655D : data <= 8'b00000000 ;
			15'h0000655E : data <= 8'b00000000 ;
			15'h0000655F : data <= 8'b00000000 ;
			15'h00006560 : data <= 8'b00000000 ;
			15'h00006561 : data <= 8'b00000000 ;
			15'h00006562 : data <= 8'b00000000 ;
			15'h00006563 : data <= 8'b00000000 ;
			15'h00006564 : data <= 8'b00000000 ;
			15'h00006565 : data <= 8'b00000000 ;
			15'h00006566 : data <= 8'b00000000 ;
			15'h00006567 : data <= 8'b00000000 ;
			15'h00006568 : data <= 8'b00000000 ;
			15'h00006569 : data <= 8'b00000000 ;
			15'h0000656A : data <= 8'b00000000 ;
			15'h0000656B : data <= 8'b00000000 ;
			15'h0000656C : data <= 8'b00000000 ;
			15'h0000656D : data <= 8'b00000000 ;
			15'h0000656E : data <= 8'b00000000 ;
			15'h0000656F : data <= 8'b00000000 ;
			15'h00006570 : data <= 8'b00000000 ;
			15'h00006571 : data <= 8'b00000000 ;
			15'h00006572 : data <= 8'b00000000 ;
			15'h00006573 : data <= 8'b00000000 ;
			15'h00006574 : data <= 8'b00000000 ;
			15'h00006575 : data <= 8'b00000000 ;
			15'h00006576 : data <= 8'b00000000 ;
			15'h00006577 : data <= 8'b00000000 ;
			15'h00006578 : data <= 8'b00000000 ;
			15'h00006579 : data <= 8'b00000000 ;
			15'h0000657A : data <= 8'b00000000 ;
			15'h0000657B : data <= 8'b00000000 ;
			15'h0000657C : data <= 8'b00000000 ;
			15'h0000657D : data <= 8'b00000000 ;
			15'h0000657E : data <= 8'b00000000 ;
			15'h0000657F : data <= 8'b00000000 ;
			15'h00006580 : data <= 8'b00000000 ;
			15'h00006581 : data <= 8'b00000000 ;
			15'h00006582 : data <= 8'b00000000 ;
			15'h00006583 : data <= 8'b00000000 ;
			15'h00006584 : data <= 8'b00000000 ;
			15'h00006585 : data <= 8'b00000000 ;
			15'h00006586 : data <= 8'b00000000 ;
			15'h00006587 : data <= 8'b00000000 ;
			15'h00006588 : data <= 8'b00000000 ;
			15'h00006589 : data <= 8'b00000000 ;
			15'h0000658A : data <= 8'b00000000 ;
			15'h0000658B : data <= 8'b00000000 ;
			15'h0000658C : data <= 8'b00000000 ;
			15'h0000658D : data <= 8'b00000000 ;
			15'h0000658E : data <= 8'b00000000 ;
			15'h0000658F : data <= 8'b00000000 ;
			15'h00006590 : data <= 8'b00000000 ;
			15'h00006591 : data <= 8'b00000000 ;
			15'h00006592 : data <= 8'b00000000 ;
			15'h00006593 : data <= 8'b00000000 ;
			15'h00006594 : data <= 8'b00000000 ;
			15'h00006595 : data <= 8'b00000000 ;
			15'h00006596 : data <= 8'b00000000 ;
			15'h00006597 : data <= 8'b00000000 ;
			15'h00006598 : data <= 8'b00000000 ;
			15'h00006599 : data <= 8'b00000000 ;
			15'h0000659A : data <= 8'b00000000 ;
			15'h0000659B : data <= 8'b00000000 ;
			15'h0000659C : data <= 8'b00000000 ;
			15'h0000659D : data <= 8'b00000000 ;
			15'h0000659E : data <= 8'b00000000 ;
			15'h0000659F : data <= 8'b00000000 ;
			15'h000065A0 : data <= 8'b00000000 ;
			15'h000065A1 : data <= 8'b00000000 ;
			15'h000065A2 : data <= 8'b00000000 ;
			15'h000065A3 : data <= 8'b00000000 ;
			15'h000065A4 : data <= 8'b00000000 ;
			15'h000065A5 : data <= 8'b00000000 ;
			15'h000065A6 : data <= 8'b00000000 ;
			15'h000065A7 : data <= 8'b00000000 ;
			15'h000065A8 : data <= 8'b00000000 ;
			15'h000065A9 : data <= 8'b00000000 ;
			15'h000065AA : data <= 8'b00000000 ;
			15'h000065AB : data <= 8'b00000000 ;
			15'h000065AC : data <= 8'b00000000 ;
			15'h000065AD : data <= 8'b00000000 ;
			15'h000065AE : data <= 8'b00000000 ;
			15'h000065AF : data <= 8'b00000000 ;
			15'h000065B0 : data <= 8'b00000000 ;
			15'h000065B1 : data <= 8'b00000000 ;
			15'h000065B2 : data <= 8'b00000000 ;
			15'h000065B3 : data <= 8'b00000000 ;
			15'h000065B4 : data <= 8'b00000000 ;
			15'h000065B5 : data <= 8'b00000000 ;
			15'h000065B6 : data <= 8'b00000000 ;
			15'h000065B7 : data <= 8'b00000000 ;
			15'h000065B8 : data <= 8'b00000000 ;
			15'h000065B9 : data <= 8'b00000000 ;
			15'h000065BA : data <= 8'b00000000 ;
			15'h000065BB : data <= 8'b00000000 ;
			15'h000065BC : data <= 8'b00000000 ;
			15'h000065BD : data <= 8'b00000000 ;
			15'h000065BE : data <= 8'b00000000 ;
			15'h000065BF : data <= 8'b00000000 ;
			15'h000065C0 : data <= 8'b00000000 ;
			15'h000065C1 : data <= 8'b00000000 ;
			15'h000065C2 : data <= 8'b00000000 ;
			15'h000065C3 : data <= 8'b00000000 ;
			15'h000065C4 : data <= 8'b00000000 ;
			15'h000065C5 : data <= 8'b00000000 ;
			15'h000065C6 : data <= 8'b00000000 ;
			15'h000065C7 : data <= 8'b00000000 ;
			15'h000065C8 : data <= 8'b00000000 ;
			15'h000065C9 : data <= 8'b00000000 ;
			15'h000065CA : data <= 8'b00000000 ;
			15'h000065CB : data <= 8'b00000000 ;
			15'h000065CC : data <= 8'b00000000 ;
			15'h000065CD : data <= 8'b00000000 ;
			15'h000065CE : data <= 8'b00000000 ;
			15'h000065CF : data <= 8'b00000000 ;
			15'h000065D0 : data <= 8'b00000000 ;
			15'h000065D1 : data <= 8'b00000000 ;
			15'h000065D2 : data <= 8'b00000000 ;
			15'h000065D3 : data <= 8'b00000000 ;
			15'h000065D4 : data <= 8'b00000000 ;
			15'h000065D5 : data <= 8'b00000000 ;
			15'h000065D6 : data <= 8'b00000000 ;
			15'h000065D7 : data <= 8'b00000000 ;
			15'h000065D8 : data <= 8'b00000000 ;
			15'h000065D9 : data <= 8'b00000000 ;
			15'h000065DA : data <= 8'b00000000 ;
			15'h000065DB : data <= 8'b00000000 ;
			15'h000065DC : data <= 8'b00000000 ;
			15'h000065DD : data <= 8'b00000000 ;
			15'h000065DE : data <= 8'b00000000 ;
			15'h000065DF : data <= 8'b00000000 ;
			15'h000065E0 : data <= 8'b00000000 ;
			15'h000065E1 : data <= 8'b00000000 ;
			15'h000065E2 : data <= 8'b00000000 ;
			15'h000065E3 : data <= 8'b00000000 ;
			15'h000065E4 : data <= 8'b00000000 ;
			15'h000065E5 : data <= 8'b00000000 ;
			15'h000065E6 : data <= 8'b00000000 ;
			15'h000065E7 : data <= 8'b00000000 ;
			15'h000065E8 : data <= 8'b00000000 ;
			15'h000065E9 : data <= 8'b00000000 ;
			15'h000065EA : data <= 8'b00000000 ;
			15'h000065EB : data <= 8'b00000000 ;
			15'h000065EC : data <= 8'b00000000 ;
			15'h000065ED : data <= 8'b00000000 ;
			15'h000065EE : data <= 8'b00000000 ;
			15'h000065EF : data <= 8'b00000000 ;
			15'h000065F0 : data <= 8'b00000000 ;
			15'h000065F1 : data <= 8'b00000000 ;
			15'h000065F2 : data <= 8'b00000000 ;
			15'h000065F3 : data <= 8'b00000000 ;
			15'h000065F4 : data <= 8'b00000000 ;
			15'h000065F5 : data <= 8'b00000000 ;
			15'h000065F6 : data <= 8'b00000000 ;
			15'h000065F7 : data <= 8'b00000000 ;
			15'h000065F8 : data <= 8'b00000000 ;
			15'h000065F9 : data <= 8'b00000000 ;
			15'h000065FA : data <= 8'b00000000 ;
			15'h000065FB : data <= 8'b00000000 ;
			15'h000065FC : data <= 8'b00000000 ;
			15'h000065FD : data <= 8'b00000000 ;
			15'h000065FE : data <= 8'b00000000 ;
			15'h000065FF : data <= 8'b00000000 ;
			15'h00006600 : data <= 8'b00000000 ;
			15'h00006601 : data <= 8'b00000000 ;
			15'h00006602 : data <= 8'b00000000 ;
			15'h00006603 : data <= 8'b00000000 ;
			15'h00006604 : data <= 8'b00000000 ;
			15'h00006605 : data <= 8'b00000000 ;
			15'h00006606 : data <= 8'b00000000 ;
			15'h00006607 : data <= 8'b00000000 ;
			15'h00006608 : data <= 8'b00000000 ;
			15'h00006609 : data <= 8'b00000000 ;
			15'h0000660A : data <= 8'b00000000 ;
			15'h0000660B : data <= 8'b00000000 ;
			15'h0000660C : data <= 8'b00000000 ;
			15'h0000660D : data <= 8'b00000000 ;
			15'h0000660E : data <= 8'b00000000 ;
			15'h0000660F : data <= 8'b00000000 ;
			15'h00006610 : data <= 8'b00000000 ;
			15'h00006611 : data <= 8'b00000000 ;
			15'h00006612 : data <= 8'b00000000 ;
			15'h00006613 : data <= 8'b00000000 ;
			15'h00006614 : data <= 8'b00000000 ;
			15'h00006615 : data <= 8'b00000000 ;
			15'h00006616 : data <= 8'b00000000 ;
			15'h00006617 : data <= 8'b00000000 ;
			15'h00006618 : data <= 8'b00000000 ;
			15'h00006619 : data <= 8'b00000000 ;
			15'h0000661A : data <= 8'b00000000 ;
			15'h0000661B : data <= 8'b00000000 ;
			15'h0000661C : data <= 8'b00000000 ;
			15'h0000661D : data <= 8'b00000000 ;
			15'h0000661E : data <= 8'b00000000 ;
			15'h0000661F : data <= 8'b00000000 ;
			15'h00006620 : data <= 8'b00000000 ;
			15'h00006621 : data <= 8'b00000000 ;
			15'h00006622 : data <= 8'b00000000 ;
			15'h00006623 : data <= 8'b00000000 ;
			15'h00006624 : data <= 8'b00000000 ;
			15'h00006625 : data <= 8'b00000000 ;
			15'h00006626 : data <= 8'b00000000 ;
			15'h00006627 : data <= 8'b00000000 ;
			15'h00006628 : data <= 8'b00000000 ;
			15'h00006629 : data <= 8'b00000000 ;
			15'h0000662A : data <= 8'b00000000 ;
			15'h0000662B : data <= 8'b00000000 ;
			15'h0000662C : data <= 8'b00000000 ;
			15'h0000662D : data <= 8'b00000000 ;
			15'h0000662E : data <= 8'b00000000 ;
			15'h0000662F : data <= 8'b00000000 ;
			15'h00006630 : data <= 8'b00000000 ;
			15'h00006631 : data <= 8'b00000000 ;
			15'h00006632 : data <= 8'b00000000 ;
			15'h00006633 : data <= 8'b00000000 ;
			15'h00006634 : data <= 8'b00000000 ;
			15'h00006635 : data <= 8'b00000000 ;
			15'h00006636 : data <= 8'b00000000 ;
			15'h00006637 : data <= 8'b00000000 ;
			15'h00006638 : data <= 8'b00000000 ;
			15'h00006639 : data <= 8'b00000000 ;
			15'h0000663A : data <= 8'b00000000 ;
			15'h0000663B : data <= 8'b00000000 ;
			15'h0000663C : data <= 8'b00000000 ;
			15'h0000663D : data <= 8'b00000000 ;
			15'h0000663E : data <= 8'b00000000 ;
			15'h0000663F : data <= 8'b00000000 ;
			15'h00006640 : data <= 8'b00000000 ;
			15'h00006641 : data <= 8'b00000000 ;
			15'h00006642 : data <= 8'b00000000 ;
			15'h00006643 : data <= 8'b00000000 ;
			15'h00006644 : data <= 8'b00000000 ;
			15'h00006645 : data <= 8'b00000000 ;
			15'h00006646 : data <= 8'b00000000 ;
			15'h00006647 : data <= 8'b00000000 ;
			15'h00006648 : data <= 8'b00000000 ;
			15'h00006649 : data <= 8'b00000000 ;
			15'h0000664A : data <= 8'b00000000 ;
			15'h0000664B : data <= 8'b00000000 ;
			15'h0000664C : data <= 8'b00000000 ;
			15'h0000664D : data <= 8'b00000000 ;
			15'h0000664E : data <= 8'b00000000 ;
			15'h0000664F : data <= 8'b00000000 ;
			15'h00006650 : data <= 8'b00000000 ;
			15'h00006651 : data <= 8'b00000000 ;
			15'h00006652 : data <= 8'b00000000 ;
			15'h00006653 : data <= 8'b00000000 ;
			15'h00006654 : data <= 8'b00000000 ;
			15'h00006655 : data <= 8'b00000000 ;
			15'h00006656 : data <= 8'b00000000 ;
			15'h00006657 : data <= 8'b00000000 ;
			15'h00006658 : data <= 8'b00000000 ;
			15'h00006659 : data <= 8'b00000000 ;
			15'h0000665A : data <= 8'b00000000 ;
			15'h0000665B : data <= 8'b00000000 ;
			15'h0000665C : data <= 8'b00000000 ;
			15'h0000665D : data <= 8'b00000000 ;
			15'h0000665E : data <= 8'b00000000 ;
			15'h0000665F : data <= 8'b00000000 ;
			15'h00006660 : data <= 8'b00000000 ;
			15'h00006661 : data <= 8'b00000000 ;
			15'h00006662 : data <= 8'b00000000 ;
			15'h00006663 : data <= 8'b00000000 ;
			15'h00006664 : data <= 8'b00000000 ;
			15'h00006665 : data <= 8'b00000000 ;
			15'h00006666 : data <= 8'b00000000 ;
			15'h00006667 : data <= 8'b00000000 ;
			15'h00006668 : data <= 8'b00000000 ;
			15'h00006669 : data <= 8'b00000000 ;
			15'h0000666A : data <= 8'b00000000 ;
			15'h0000666B : data <= 8'b00000000 ;
			15'h0000666C : data <= 8'b00000000 ;
			15'h0000666D : data <= 8'b00000000 ;
			15'h0000666E : data <= 8'b00000000 ;
			15'h0000666F : data <= 8'b00000000 ;
			15'h00006670 : data <= 8'b00000000 ;
			15'h00006671 : data <= 8'b00000000 ;
			15'h00006672 : data <= 8'b00000000 ;
			15'h00006673 : data <= 8'b00000000 ;
			15'h00006674 : data <= 8'b00000000 ;
			15'h00006675 : data <= 8'b00000000 ;
			15'h00006676 : data <= 8'b00000000 ;
			15'h00006677 : data <= 8'b00000000 ;
			15'h00006678 : data <= 8'b00000000 ;
			15'h00006679 : data <= 8'b00000000 ;
			15'h0000667A : data <= 8'b00000000 ;
			15'h0000667B : data <= 8'b00000000 ;
			15'h0000667C : data <= 8'b00000000 ;
			15'h0000667D : data <= 8'b00000000 ;
			15'h0000667E : data <= 8'b00000000 ;
			15'h0000667F : data <= 8'b00000000 ;
			15'h00006680 : data <= 8'b00000000 ;
			15'h00006681 : data <= 8'b00000000 ;
			15'h00006682 : data <= 8'b00000000 ;
			15'h00006683 : data <= 8'b00000000 ;
			15'h00006684 : data <= 8'b00000000 ;
			15'h00006685 : data <= 8'b00000000 ;
			15'h00006686 : data <= 8'b00000000 ;
			15'h00006687 : data <= 8'b00000000 ;
			15'h00006688 : data <= 8'b00000000 ;
			15'h00006689 : data <= 8'b00000000 ;
			15'h0000668A : data <= 8'b00000000 ;
			15'h0000668B : data <= 8'b00000000 ;
			15'h0000668C : data <= 8'b00000000 ;
			15'h0000668D : data <= 8'b00000000 ;
			15'h0000668E : data <= 8'b00000000 ;
			15'h0000668F : data <= 8'b00000000 ;
			15'h00006690 : data <= 8'b00000000 ;
			15'h00006691 : data <= 8'b00000000 ;
			15'h00006692 : data <= 8'b00000000 ;
			15'h00006693 : data <= 8'b00000000 ;
			15'h00006694 : data <= 8'b00000000 ;
			15'h00006695 : data <= 8'b00000000 ;
			15'h00006696 : data <= 8'b00000000 ;
			15'h00006697 : data <= 8'b00000000 ;
			15'h00006698 : data <= 8'b00000000 ;
			15'h00006699 : data <= 8'b00000000 ;
			15'h0000669A : data <= 8'b00000000 ;
			15'h0000669B : data <= 8'b00000000 ;
			15'h0000669C : data <= 8'b00000000 ;
			15'h0000669D : data <= 8'b00000000 ;
			15'h0000669E : data <= 8'b00000000 ;
			15'h0000669F : data <= 8'b00000000 ;
			15'h000066A0 : data <= 8'b00000000 ;
			15'h000066A1 : data <= 8'b00000000 ;
			15'h000066A2 : data <= 8'b00000000 ;
			15'h000066A3 : data <= 8'b00000000 ;
			15'h000066A4 : data <= 8'b00000000 ;
			15'h000066A5 : data <= 8'b00000000 ;
			15'h000066A6 : data <= 8'b00000000 ;
			15'h000066A7 : data <= 8'b00000000 ;
			15'h000066A8 : data <= 8'b00000000 ;
			15'h000066A9 : data <= 8'b00000000 ;
			15'h000066AA : data <= 8'b00000000 ;
			15'h000066AB : data <= 8'b00000000 ;
			15'h000066AC : data <= 8'b00000000 ;
			15'h000066AD : data <= 8'b00000000 ;
			15'h000066AE : data <= 8'b00000000 ;
			15'h000066AF : data <= 8'b00000000 ;
			15'h000066B0 : data <= 8'b00000000 ;
			15'h000066B1 : data <= 8'b00000000 ;
			15'h000066B2 : data <= 8'b00000000 ;
			15'h000066B3 : data <= 8'b00000000 ;
			15'h000066B4 : data <= 8'b00000000 ;
			15'h000066B5 : data <= 8'b00000000 ;
			15'h000066B6 : data <= 8'b00000000 ;
			15'h000066B7 : data <= 8'b00000000 ;
			15'h000066B8 : data <= 8'b00000000 ;
			15'h000066B9 : data <= 8'b00000000 ;
			15'h000066BA : data <= 8'b00000000 ;
			15'h000066BB : data <= 8'b00000000 ;
			15'h000066BC : data <= 8'b00000000 ;
			15'h000066BD : data <= 8'b00000000 ;
			15'h000066BE : data <= 8'b00000000 ;
			15'h000066BF : data <= 8'b00000000 ;
			15'h000066C0 : data <= 8'b00000000 ;
			15'h000066C1 : data <= 8'b00000000 ;
			15'h000066C2 : data <= 8'b00000000 ;
			15'h000066C3 : data <= 8'b00000000 ;
			15'h000066C4 : data <= 8'b00000000 ;
			15'h000066C5 : data <= 8'b00000000 ;
			15'h000066C6 : data <= 8'b00000000 ;
			15'h000066C7 : data <= 8'b00000000 ;
			15'h000066C8 : data <= 8'b00000000 ;
			15'h000066C9 : data <= 8'b00000000 ;
			15'h000066CA : data <= 8'b00000000 ;
			15'h000066CB : data <= 8'b00000000 ;
			15'h000066CC : data <= 8'b00000000 ;
			15'h000066CD : data <= 8'b00000000 ;
			15'h000066CE : data <= 8'b00000000 ;
			15'h000066CF : data <= 8'b00000000 ;
			15'h000066D0 : data <= 8'b00000000 ;
			15'h000066D1 : data <= 8'b00000000 ;
			15'h000066D2 : data <= 8'b00000000 ;
			15'h000066D3 : data <= 8'b00000000 ;
			15'h000066D4 : data <= 8'b00000000 ;
			15'h000066D5 : data <= 8'b00000000 ;
			15'h000066D6 : data <= 8'b00000000 ;
			15'h000066D7 : data <= 8'b00000000 ;
			15'h000066D8 : data <= 8'b00000000 ;
			15'h000066D9 : data <= 8'b00000000 ;
			15'h000066DA : data <= 8'b00000000 ;
			15'h000066DB : data <= 8'b00000000 ;
			15'h000066DC : data <= 8'b00000000 ;
			15'h000066DD : data <= 8'b00000000 ;
			15'h000066DE : data <= 8'b00000000 ;
			15'h000066DF : data <= 8'b00000000 ;
			15'h000066E0 : data <= 8'b00000000 ;
			15'h000066E1 : data <= 8'b00000000 ;
			15'h000066E2 : data <= 8'b00000000 ;
			15'h000066E3 : data <= 8'b00000000 ;
			15'h000066E4 : data <= 8'b00000000 ;
			15'h000066E5 : data <= 8'b00000000 ;
			15'h000066E6 : data <= 8'b00000000 ;
			15'h000066E7 : data <= 8'b00000000 ;
			15'h000066E8 : data <= 8'b00000000 ;
			15'h000066E9 : data <= 8'b00000000 ;
			15'h000066EA : data <= 8'b00000000 ;
			15'h000066EB : data <= 8'b00000000 ;
			15'h000066EC : data <= 8'b00000000 ;
			15'h000066ED : data <= 8'b00000000 ;
			15'h000066EE : data <= 8'b00000000 ;
			15'h000066EF : data <= 8'b00000000 ;
			15'h000066F0 : data <= 8'b00000000 ;
			15'h000066F1 : data <= 8'b00000000 ;
			15'h000066F2 : data <= 8'b00000000 ;
			15'h000066F3 : data <= 8'b00000000 ;
			15'h000066F4 : data <= 8'b00000000 ;
			15'h000066F5 : data <= 8'b00000000 ;
			15'h000066F6 : data <= 8'b00000000 ;
			15'h000066F7 : data <= 8'b00000000 ;
			15'h000066F8 : data <= 8'b00000000 ;
			15'h000066F9 : data <= 8'b00000000 ;
			15'h000066FA : data <= 8'b00000000 ;
			15'h000066FB : data <= 8'b00000000 ;
			15'h000066FC : data <= 8'b00000000 ;
			15'h000066FD : data <= 8'b00000000 ;
			15'h000066FE : data <= 8'b00000000 ;
			15'h000066FF : data <= 8'b00000000 ;
			15'h00006700 : data <= 8'b00000000 ;
			15'h00006701 : data <= 8'b00000000 ;
			15'h00006702 : data <= 8'b00000000 ;
			15'h00006703 : data <= 8'b00000000 ;
			15'h00006704 : data <= 8'b00000000 ;
			15'h00006705 : data <= 8'b00000000 ;
			15'h00006706 : data <= 8'b00000000 ;
			15'h00006707 : data <= 8'b00000000 ;
			15'h00006708 : data <= 8'b00000000 ;
			15'h00006709 : data <= 8'b00000000 ;
			15'h0000670A : data <= 8'b00000000 ;
			15'h0000670B : data <= 8'b00000000 ;
			15'h0000670C : data <= 8'b00000000 ;
			15'h0000670D : data <= 8'b00000000 ;
			15'h0000670E : data <= 8'b00000000 ;
			15'h0000670F : data <= 8'b00000000 ;
			15'h00006710 : data <= 8'b00000000 ;
			15'h00006711 : data <= 8'b00000000 ;
			15'h00006712 : data <= 8'b00000000 ;
			15'h00006713 : data <= 8'b00000000 ;
			15'h00006714 : data <= 8'b00000000 ;
			15'h00006715 : data <= 8'b00000000 ;
			15'h00006716 : data <= 8'b00000000 ;
			15'h00006717 : data <= 8'b00000000 ;
			15'h00006718 : data <= 8'b00000000 ;
			15'h00006719 : data <= 8'b00000000 ;
			15'h0000671A : data <= 8'b00000000 ;
			15'h0000671B : data <= 8'b00000000 ;
			15'h0000671C : data <= 8'b00000000 ;
			15'h0000671D : data <= 8'b00000000 ;
			15'h0000671E : data <= 8'b00000000 ;
			15'h0000671F : data <= 8'b00000000 ;
			15'h00006720 : data <= 8'b00000000 ;
			15'h00006721 : data <= 8'b00000000 ;
			15'h00006722 : data <= 8'b00000000 ;
			15'h00006723 : data <= 8'b00000000 ;
			15'h00006724 : data <= 8'b00000000 ;
			15'h00006725 : data <= 8'b00000000 ;
			15'h00006726 : data <= 8'b00000000 ;
			15'h00006727 : data <= 8'b00000000 ;
			15'h00006728 : data <= 8'b00000000 ;
			15'h00006729 : data <= 8'b00000000 ;
			15'h0000672A : data <= 8'b00000000 ;
			15'h0000672B : data <= 8'b00000000 ;
			15'h0000672C : data <= 8'b00000000 ;
			15'h0000672D : data <= 8'b00000000 ;
			15'h0000672E : data <= 8'b00000000 ;
			15'h0000672F : data <= 8'b00000000 ;
			15'h00006730 : data <= 8'b00000000 ;
			15'h00006731 : data <= 8'b00000000 ;
			15'h00006732 : data <= 8'b00000000 ;
			15'h00006733 : data <= 8'b00000000 ;
			15'h00006734 : data <= 8'b00000000 ;
			15'h00006735 : data <= 8'b00000000 ;
			15'h00006736 : data <= 8'b00000000 ;
			15'h00006737 : data <= 8'b00000000 ;
			15'h00006738 : data <= 8'b00000000 ;
			15'h00006739 : data <= 8'b00000000 ;
			15'h0000673A : data <= 8'b00000000 ;
			15'h0000673B : data <= 8'b00000000 ;
			15'h0000673C : data <= 8'b00000000 ;
			15'h0000673D : data <= 8'b00000000 ;
			15'h0000673E : data <= 8'b00000000 ;
			15'h0000673F : data <= 8'b00000000 ;
			15'h00006740 : data <= 8'b00000000 ;
			15'h00006741 : data <= 8'b00000000 ;
			15'h00006742 : data <= 8'b00000000 ;
			15'h00006743 : data <= 8'b00000000 ;
			15'h00006744 : data <= 8'b00000000 ;
			15'h00006745 : data <= 8'b00000000 ;
			15'h00006746 : data <= 8'b00000000 ;
			15'h00006747 : data <= 8'b00000000 ;
			15'h00006748 : data <= 8'b00000000 ;
			15'h00006749 : data <= 8'b00000000 ;
			15'h0000674A : data <= 8'b00000000 ;
			15'h0000674B : data <= 8'b00000000 ;
			15'h0000674C : data <= 8'b00000000 ;
			15'h0000674D : data <= 8'b00000000 ;
			15'h0000674E : data <= 8'b00000000 ;
			15'h0000674F : data <= 8'b00000000 ;
			15'h00006750 : data <= 8'b00000000 ;
			15'h00006751 : data <= 8'b00000000 ;
			15'h00006752 : data <= 8'b00000000 ;
			15'h00006753 : data <= 8'b00000000 ;
			15'h00006754 : data <= 8'b00000000 ;
			15'h00006755 : data <= 8'b00000000 ;
			15'h00006756 : data <= 8'b00000000 ;
			15'h00006757 : data <= 8'b00000000 ;
			15'h00006758 : data <= 8'b00000000 ;
			15'h00006759 : data <= 8'b00000000 ;
			15'h0000675A : data <= 8'b00000000 ;
			15'h0000675B : data <= 8'b00000000 ;
			15'h0000675C : data <= 8'b00000000 ;
			15'h0000675D : data <= 8'b00000000 ;
			15'h0000675E : data <= 8'b00000000 ;
			15'h0000675F : data <= 8'b00000000 ;
			15'h00006760 : data <= 8'b00000000 ;
			15'h00006761 : data <= 8'b00000000 ;
			15'h00006762 : data <= 8'b00000000 ;
			15'h00006763 : data <= 8'b00000000 ;
			15'h00006764 : data <= 8'b00000000 ;
			15'h00006765 : data <= 8'b00000000 ;
			15'h00006766 : data <= 8'b00000000 ;
			15'h00006767 : data <= 8'b00000000 ;
			15'h00006768 : data <= 8'b00000000 ;
			15'h00006769 : data <= 8'b00000000 ;
			15'h0000676A : data <= 8'b00000000 ;
			15'h0000676B : data <= 8'b00000000 ;
			15'h0000676C : data <= 8'b00000000 ;
			15'h0000676D : data <= 8'b00000000 ;
			15'h0000676E : data <= 8'b00000000 ;
			15'h0000676F : data <= 8'b00000000 ;
			15'h00006770 : data <= 8'b00000000 ;
			15'h00006771 : data <= 8'b00000000 ;
			15'h00006772 : data <= 8'b00000000 ;
			15'h00006773 : data <= 8'b00000000 ;
			15'h00006774 : data <= 8'b00000000 ;
			15'h00006775 : data <= 8'b00000000 ;
			15'h00006776 : data <= 8'b00000000 ;
			15'h00006777 : data <= 8'b00000000 ;
			15'h00006778 : data <= 8'b00000000 ;
			15'h00006779 : data <= 8'b00000000 ;
			15'h0000677A : data <= 8'b00000000 ;
			15'h0000677B : data <= 8'b00000000 ;
			15'h0000677C : data <= 8'b00000000 ;
			15'h0000677D : data <= 8'b00000000 ;
			15'h0000677E : data <= 8'b00000000 ;
			15'h0000677F : data <= 8'b00000000 ;
			15'h00006780 : data <= 8'b00000000 ;
			15'h00006781 : data <= 8'b00000000 ;
			15'h00006782 : data <= 8'b00000000 ;
			15'h00006783 : data <= 8'b00000000 ;
			15'h00006784 : data <= 8'b00000000 ;
			15'h00006785 : data <= 8'b00000000 ;
			15'h00006786 : data <= 8'b00000000 ;
			15'h00006787 : data <= 8'b00000000 ;
			15'h00006788 : data <= 8'b00000000 ;
			15'h00006789 : data <= 8'b00000000 ;
			15'h0000678A : data <= 8'b00000000 ;
			15'h0000678B : data <= 8'b00000000 ;
			15'h0000678C : data <= 8'b00000000 ;
			15'h0000678D : data <= 8'b00000000 ;
			15'h0000678E : data <= 8'b00000000 ;
			15'h0000678F : data <= 8'b00000000 ;
			15'h00006790 : data <= 8'b00000000 ;
			15'h00006791 : data <= 8'b00000000 ;
			15'h00006792 : data <= 8'b00000000 ;
			15'h00006793 : data <= 8'b00000000 ;
			15'h00006794 : data <= 8'b00000000 ;
			15'h00006795 : data <= 8'b00000000 ;
			15'h00006796 : data <= 8'b00000000 ;
			15'h00006797 : data <= 8'b00000000 ;
			15'h00006798 : data <= 8'b00000000 ;
			15'h00006799 : data <= 8'b00000000 ;
			15'h0000679A : data <= 8'b00000000 ;
			15'h0000679B : data <= 8'b00000000 ;
			15'h0000679C : data <= 8'b00000000 ;
			15'h0000679D : data <= 8'b00000000 ;
			15'h0000679E : data <= 8'b00000000 ;
			15'h0000679F : data <= 8'b00000000 ;
			15'h000067A0 : data <= 8'b00000000 ;
			15'h000067A1 : data <= 8'b00000000 ;
			15'h000067A2 : data <= 8'b00000000 ;
			15'h000067A3 : data <= 8'b00000000 ;
			15'h000067A4 : data <= 8'b00000000 ;
			15'h000067A5 : data <= 8'b00000000 ;
			15'h000067A6 : data <= 8'b00000000 ;
			15'h000067A7 : data <= 8'b00000000 ;
			15'h000067A8 : data <= 8'b00000000 ;
			15'h000067A9 : data <= 8'b00000000 ;
			15'h000067AA : data <= 8'b00000000 ;
			15'h000067AB : data <= 8'b00000000 ;
			15'h000067AC : data <= 8'b00000000 ;
			15'h000067AD : data <= 8'b00000000 ;
			15'h000067AE : data <= 8'b00000000 ;
			15'h000067AF : data <= 8'b00000000 ;
			15'h000067B0 : data <= 8'b00000000 ;
			15'h000067B1 : data <= 8'b00000000 ;
			15'h000067B2 : data <= 8'b00000000 ;
			15'h000067B3 : data <= 8'b00000000 ;
			15'h000067B4 : data <= 8'b00000000 ;
			15'h000067B5 : data <= 8'b00000000 ;
			15'h000067B6 : data <= 8'b00000000 ;
			15'h000067B7 : data <= 8'b00000000 ;
			15'h000067B8 : data <= 8'b00000000 ;
			15'h000067B9 : data <= 8'b00000000 ;
			15'h000067BA : data <= 8'b00000000 ;
			15'h000067BB : data <= 8'b00000000 ;
			15'h000067BC : data <= 8'b00000000 ;
			15'h000067BD : data <= 8'b00000000 ;
			15'h000067BE : data <= 8'b00000000 ;
			15'h000067BF : data <= 8'b00000000 ;
			15'h000067C0 : data <= 8'b00000000 ;
			15'h000067C1 : data <= 8'b00000000 ;
			15'h000067C2 : data <= 8'b00000000 ;
			15'h000067C3 : data <= 8'b00000000 ;
			15'h000067C4 : data <= 8'b00000000 ;
			15'h000067C5 : data <= 8'b00000000 ;
			15'h000067C6 : data <= 8'b00000000 ;
			15'h000067C7 : data <= 8'b00000000 ;
			15'h000067C8 : data <= 8'b00000000 ;
			15'h000067C9 : data <= 8'b00000000 ;
			15'h000067CA : data <= 8'b00000000 ;
			15'h000067CB : data <= 8'b00000000 ;
			15'h000067CC : data <= 8'b00000000 ;
			15'h000067CD : data <= 8'b00000000 ;
			15'h000067CE : data <= 8'b00000000 ;
			15'h000067CF : data <= 8'b00000000 ;
			15'h000067D0 : data <= 8'b00000000 ;
			15'h000067D1 : data <= 8'b00000000 ;
			15'h000067D2 : data <= 8'b00000000 ;
			15'h000067D3 : data <= 8'b00000000 ;
			15'h000067D4 : data <= 8'b00000000 ;
			15'h000067D5 : data <= 8'b00000000 ;
			15'h000067D6 : data <= 8'b00000000 ;
			15'h000067D7 : data <= 8'b00000000 ;
			15'h000067D8 : data <= 8'b00000000 ;
			15'h000067D9 : data <= 8'b00000000 ;
			15'h000067DA : data <= 8'b00000000 ;
			15'h000067DB : data <= 8'b00000000 ;
			15'h000067DC : data <= 8'b00000000 ;
			15'h000067DD : data <= 8'b00000000 ;
			15'h000067DE : data <= 8'b00000000 ;
			15'h000067DF : data <= 8'b00000000 ;
			15'h000067E0 : data <= 8'b00000000 ;
			15'h000067E1 : data <= 8'b00000000 ;
			15'h000067E2 : data <= 8'b00000000 ;
			15'h000067E3 : data <= 8'b00000000 ;
			15'h000067E4 : data <= 8'b00000000 ;
			15'h000067E5 : data <= 8'b00000000 ;
			15'h000067E6 : data <= 8'b00000000 ;
			15'h000067E7 : data <= 8'b00000000 ;
			15'h000067E8 : data <= 8'b00000000 ;
			15'h000067E9 : data <= 8'b00000000 ;
			15'h000067EA : data <= 8'b00000000 ;
			15'h000067EB : data <= 8'b00000000 ;
			15'h000067EC : data <= 8'b00000000 ;
			15'h000067ED : data <= 8'b00000000 ;
			15'h000067EE : data <= 8'b00000000 ;
			15'h000067EF : data <= 8'b00000000 ;
			15'h000067F0 : data <= 8'b00000000 ;
			15'h000067F1 : data <= 8'b00000000 ;
			15'h000067F2 : data <= 8'b00000000 ;
			15'h000067F3 : data <= 8'b00000000 ;
			15'h000067F4 : data <= 8'b00000000 ;
			15'h000067F5 : data <= 8'b00000000 ;
			15'h000067F6 : data <= 8'b00000000 ;
			15'h000067F7 : data <= 8'b00000000 ;
			15'h000067F8 : data <= 8'b00000000 ;
			15'h000067F9 : data <= 8'b00000000 ;
			15'h000067FA : data <= 8'b00000000 ;
			15'h000067FB : data <= 8'b00000000 ;
			15'h000067FC : data <= 8'b00000000 ;
			15'h000067FD : data <= 8'b00000000 ;
			15'h000067FE : data <= 8'b00000000 ;
			15'h000067FF : data <= 8'b00000000 ;
			15'h00006800 : data <= 8'b00000000 ;
			15'h00006801 : data <= 8'b00000000 ;
			15'h00006802 : data <= 8'b00000000 ;
			15'h00006803 : data <= 8'b00000000 ;
			15'h00006804 : data <= 8'b00000000 ;
			15'h00006805 : data <= 8'b00000000 ;
			15'h00006806 : data <= 8'b00000000 ;
			15'h00006807 : data <= 8'b00000000 ;
			15'h00006808 : data <= 8'b00000000 ;
			15'h00006809 : data <= 8'b00000000 ;
			15'h0000680A : data <= 8'b00000000 ;
			15'h0000680B : data <= 8'b00000000 ;
			15'h0000680C : data <= 8'b00000000 ;
			15'h0000680D : data <= 8'b00000000 ;
			15'h0000680E : data <= 8'b00000000 ;
			15'h0000680F : data <= 8'b00000000 ;
			15'h00006810 : data <= 8'b00000000 ;
			15'h00006811 : data <= 8'b00000000 ;
			15'h00006812 : data <= 8'b00000000 ;
			15'h00006813 : data <= 8'b00000000 ;
			15'h00006814 : data <= 8'b00000000 ;
			15'h00006815 : data <= 8'b00000000 ;
			15'h00006816 : data <= 8'b00000000 ;
			15'h00006817 : data <= 8'b00000000 ;
			15'h00006818 : data <= 8'b00000000 ;
			15'h00006819 : data <= 8'b00000000 ;
			15'h0000681A : data <= 8'b00000000 ;
			15'h0000681B : data <= 8'b00000000 ;
			15'h0000681C : data <= 8'b00000000 ;
			15'h0000681D : data <= 8'b00000000 ;
			15'h0000681E : data <= 8'b00000000 ;
			15'h0000681F : data <= 8'b00000000 ;
			15'h00006820 : data <= 8'b00000000 ;
			15'h00006821 : data <= 8'b00000000 ;
			15'h00006822 : data <= 8'b00000000 ;
			15'h00006823 : data <= 8'b00000000 ;
			15'h00006824 : data <= 8'b00000000 ;
			15'h00006825 : data <= 8'b00000000 ;
			15'h00006826 : data <= 8'b00000000 ;
			15'h00006827 : data <= 8'b00000000 ;
			15'h00006828 : data <= 8'b00000000 ;
			15'h00006829 : data <= 8'b00000000 ;
			15'h0000682A : data <= 8'b00000000 ;
			15'h0000682B : data <= 8'b00000000 ;
			15'h0000682C : data <= 8'b00000000 ;
			15'h0000682D : data <= 8'b00000000 ;
			15'h0000682E : data <= 8'b00000000 ;
			15'h0000682F : data <= 8'b00000000 ;
			15'h00006830 : data <= 8'b00000000 ;
			15'h00006831 : data <= 8'b00000000 ;
			15'h00006832 : data <= 8'b00000000 ;
			15'h00006833 : data <= 8'b00000000 ;
			15'h00006834 : data <= 8'b00000000 ;
			15'h00006835 : data <= 8'b00000000 ;
			15'h00006836 : data <= 8'b00000000 ;
			15'h00006837 : data <= 8'b00000000 ;
			15'h00006838 : data <= 8'b00000000 ;
			15'h00006839 : data <= 8'b00000000 ;
			15'h0000683A : data <= 8'b00000000 ;
			15'h0000683B : data <= 8'b00000000 ;
			15'h0000683C : data <= 8'b00000000 ;
			15'h0000683D : data <= 8'b00000000 ;
			15'h0000683E : data <= 8'b00000000 ;
			15'h0000683F : data <= 8'b00000000 ;
			15'h00006840 : data <= 8'b00000000 ;
			15'h00006841 : data <= 8'b00000000 ;
			15'h00006842 : data <= 8'b00000000 ;
			15'h00006843 : data <= 8'b00000000 ;
			15'h00006844 : data <= 8'b00000000 ;
			15'h00006845 : data <= 8'b00000000 ;
			15'h00006846 : data <= 8'b00000000 ;
			15'h00006847 : data <= 8'b00000000 ;
			15'h00006848 : data <= 8'b00000000 ;
			15'h00006849 : data <= 8'b00000000 ;
			15'h0000684A : data <= 8'b00000000 ;
			15'h0000684B : data <= 8'b00000000 ;
			15'h0000684C : data <= 8'b00000000 ;
			15'h0000684D : data <= 8'b00000000 ;
			15'h0000684E : data <= 8'b00000000 ;
			15'h0000684F : data <= 8'b00000000 ;
			15'h00006850 : data <= 8'b00000000 ;
			15'h00006851 : data <= 8'b00000000 ;
			15'h00006852 : data <= 8'b00000000 ;
			15'h00006853 : data <= 8'b00000000 ;
			15'h00006854 : data <= 8'b00000000 ;
			15'h00006855 : data <= 8'b00000000 ;
			15'h00006856 : data <= 8'b00000000 ;
			15'h00006857 : data <= 8'b00000000 ;
			15'h00006858 : data <= 8'b00000000 ;
			15'h00006859 : data <= 8'b00000000 ;
			15'h0000685A : data <= 8'b00000000 ;
			15'h0000685B : data <= 8'b00000000 ;
			15'h0000685C : data <= 8'b00000000 ;
			15'h0000685D : data <= 8'b00000000 ;
			15'h0000685E : data <= 8'b00000000 ;
			15'h0000685F : data <= 8'b00000000 ;
			15'h00006860 : data <= 8'b00000000 ;
			15'h00006861 : data <= 8'b00000000 ;
			15'h00006862 : data <= 8'b00000000 ;
			15'h00006863 : data <= 8'b00000000 ;
			15'h00006864 : data <= 8'b00000000 ;
			15'h00006865 : data <= 8'b00000000 ;
			15'h00006866 : data <= 8'b00000000 ;
			15'h00006867 : data <= 8'b00000000 ;
			15'h00006868 : data <= 8'b00000000 ;
			15'h00006869 : data <= 8'b00000000 ;
			15'h0000686A : data <= 8'b00000000 ;
			15'h0000686B : data <= 8'b00000000 ;
			15'h0000686C : data <= 8'b00000000 ;
			15'h0000686D : data <= 8'b00000000 ;
			15'h0000686E : data <= 8'b00000000 ;
			15'h0000686F : data <= 8'b00000000 ;
			15'h00006870 : data <= 8'b00000000 ;
			15'h00006871 : data <= 8'b00000000 ;
			15'h00006872 : data <= 8'b00000000 ;
			15'h00006873 : data <= 8'b00000000 ;
			15'h00006874 : data <= 8'b00000000 ;
			15'h00006875 : data <= 8'b00000000 ;
			15'h00006876 : data <= 8'b00000000 ;
			15'h00006877 : data <= 8'b00000000 ;
			15'h00006878 : data <= 8'b00000000 ;
			15'h00006879 : data <= 8'b00000000 ;
			15'h0000687A : data <= 8'b00000000 ;
			15'h0000687B : data <= 8'b00000000 ;
			15'h0000687C : data <= 8'b00000000 ;
			15'h0000687D : data <= 8'b00000000 ;
			15'h0000687E : data <= 8'b00000000 ;
			15'h0000687F : data <= 8'b00000000 ;
			15'h00006880 : data <= 8'b00000000 ;
			15'h00006881 : data <= 8'b00000000 ;
			15'h00006882 : data <= 8'b00000000 ;
			15'h00006883 : data <= 8'b00000000 ;
			15'h00006884 : data <= 8'b00000000 ;
			15'h00006885 : data <= 8'b00000000 ;
			15'h00006886 : data <= 8'b00000000 ;
			15'h00006887 : data <= 8'b00000000 ;
			15'h00006888 : data <= 8'b00000000 ;
			15'h00006889 : data <= 8'b00000000 ;
			15'h0000688A : data <= 8'b00000000 ;
			15'h0000688B : data <= 8'b00000000 ;
			15'h0000688C : data <= 8'b00000000 ;
			15'h0000688D : data <= 8'b00000000 ;
			15'h0000688E : data <= 8'b00000000 ;
			15'h0000688F : data <= 8'b00000000 ;
			15'h00006890 : data <= 8'b00000000 ;
			15'h00006891 : data <= 8'b00000000 ;
			15'h00006892 : data <= 8'b00000000 ;
			15'h00006893 : data <= 8'b00000000 ;
			15'h00006894 : data <= 8'b00000000 ;
			15'h00006895 : data <= 8'b00000000 ;
			15'h00006896 : data <= 8'b00000000 ;
			15'h00006897 : data <= 8'b00000000 ;
			15'h00006898 : data <= 8'b00000000 ;
			15'h00006899 : data <= 8'b00000000 ;
			15'h0000689A : data <= 8'b00000000 ;
			15'h0000689B : data <= 8'b00000000 ;
			15'h0000689C : data <= 8'b00000000 ;
			15'h0000689D : data <= 8'b00000000 ;
			15'h0000689E : data <= 8'b00000000 ;
			15'h0000689F : data <= 8'b00000000 ;
			15'h000068A0 : data <= 8'b00000000 ;
			15'h000068A1 : data <= 8'b00000000 ;
			15'h000068A2 : data <= 8'b00000000 ;
			15'h000068A3 : data <= 8'b00000000 ;
			15'h000068A4 : data <= 8'b00000000 ;
			15'h000068A5 : data <= 8'b00000000 ;
			15'h000068A6 : data <= 8'b00000000 ;
			15'h000068A7 : data <= 8'b00000000 ;
			15'h000068A8 : data <= 8'b00000000 ;
			15'h000068A9 : data <= 8'b00000000 ;
			15'h000068AA : data <= 8'b00000000 ;
			15'h000068AB : data <= 8'b00000000 ;
			15'h000068AC : data <= 8'b00000000 ;
			15'h000068AD : data <= 8'b00000000 ;
			15'h000068AE : data <= 8'b00000000 ;
			15'h000068AF : data <= 8'b00000000 ;
			15'h000068B0 : data <= 8'b00000000 ;
			15'h000068B1 : data <= 8'b00000000 ;
			15'h000068B2 : data <= 8'b00000000 ;
			15'h000068B3 : data <= 8'b00000000 ;
			15'h000068B4 : data <= 8'b00000000 ;
			15'h000068B5 : data <= 8'b00000000 ;
			15'h000068B6 : data <= 8'b00000000 ;
			15'h000068B7 : data <= 8'b00000000 ;
			15'h000068B8 : data <= 8'b00000000 ;
			15'h000068B9 : data <= 8'b00000000 ;
			15'h000068BA : data <= 8'b00000000 ;
			15'h000068BB : data <= 8'b00000000 ;
			15'h000068BC : data <= 8'b00000000 ;
			15'h000068BD : data <= 8'b00000000 ;
			15'h000068BE : data <= 8'b00000000 ;
			15'h000068BF : data <= 8'b00000000 ;
			15'h000068C0 : data <= 8'b00000000 ;
			15'h000068C1 : data <= 8'b00000000 ;
			15'h000068C2 : data <= 8'b00000000 ;
			15'h000068C3 : data <= 8'b00000000 ;
			15'h000068C4 : data <= 8'b00000000 ;
			15'h000068C5 : data <= 8'b00000000 ;
			15'h000068C6 : data <= 8'b00000000 ;
			15'h000068C7 : data <= 8'b00000000 ;
			15'h000068C8 : data <= 8'b00000000 ;
			15'h000068C9 : data <= 8'b00000000 ;
			15'h000068CA : data <= 8'b00000000 ;
			15'h000068CB : data <= 8'b00000000 ;
			15'h000068CC : data <= 8'b00000000 ;
			15'h000068CD : data <= 8'b00000000 ;
			15'h000068CE : data <= 8'b00000000 ;
			15'h000068CF : data <= 8'b00000000 ;
			15'h000068D0 : data <= 8'b00000000 ;
			15'h000068D1 : data <= 8'b00000000 ;
			15'h000068D2 : data <= 8'b00000000 ;
			15'h000068D3 : data <= 8'b00000000 ;
			15'h000068D4 : data <= 8'b00000000 ;
			15'h000068D5 : data <= 8'b00000000 ;
			15'h000068D6 : data <= 8'b00000000 ;
			15'h000068D7 : data <= 8'b00000000 ;
			15'h000068D8 : data <= 8'b00000000 ;
			15'h000068D9 : data <= 8'b00000000 ;
			15'h000068DA : data <= 8'b00000000 ;
			15'h000068DB : data <= 8'b00000000 ;
			15'h000068DC : data <= 8'b00000000 ;
			15'h000068DD : data <= 8'b00000000 ;
			15'h000068DE : data <= 8'b00000000 ;
			15'h000068DF : data <= 8'b00000000 ;
			15'h000068E0 : data <= 8'b00000000 ;
			15'h000068E1 : data <= 8'b00000000 ;
			15'h000068E2 : data <= 8'b00000000 ;
			15'h000068E3 : data <= 8'b00000000 ;
			15'h000068E4 : data <= 8'b00000000 ;
			15'h000068E5 : data <= 8'b00000000 ;
			15'h000068E6 : data <= 8'b00000000 ;
			15'h000068E7 : data <= 8'b00000000 ;
			15'h000068E8 : data <= 8'b00000000 ;
			15'h000068E9 : data <= 8'b00000000 ;
			15'h000068EA : data <= 8'b00000000 ;
			15'h000068EB : data <= 8'b00000000 ;
			15'h000068EC : data <= 8'b00000000 ;
			15'h000068ED : data <= 8'b00000000 ;
			15'h000068EE : data <= 8'b00000000 ;
			15'h000068EF : data <= 8'b00000000 ;
			15'h000068F0 : data <= 8'b00000000 ;
			15'h000068F1 : data <= 8'b00000000 ;
			15'h000068F2 : data <= 8'b00000000 ;
			15'h000068F3 : data <= 8'b00000000 ;
			15'h000068F4 : data <= 8'b00000000 ;
			15'h000068F5 : data <= 8'b00000000 ;
			15'h000068F6 : data <= 8'b00000000 ;
			15'h000068F7 : data <= 8'b00000000 ;
			15'h000068F8 : data <= 8'b00000000 ;
			15'h000068F9 : data <= 8'b00000000 ;
			15'h000068FA : data <= 8'b00000000 ;
			15'h000068FB : data <= 8'b00000000 ;
			15'h000068FC : data <= 8'b00000000 ;
			15'h000068FD : data <= 8'b00000000 ;
			15'h000068FE : data <= 8'b00000000 ;
			15'h000068FF : data <= 8'b00000000 ;
			15'h00006900 : data <= 8'b00000000 ;
			15'h00006901 : data <= 8'b00000000 ;
			15'h00006902 : data <= 8'b00000000 ;
			15'h00006903 : data <= 8'b00000000 ;
			15'h00006904 : data <= 8'b00000000 ;
			15'h00006905 : data <= 8'b00000000 ;
			15'h00006906 : data <= 8'b00000000 ;
			15'h00006907 : data <= 8'b00000000 ;
			15'h00006908 : data <= 8'b00000000 ;
			15'h00006909 : data <= 8'b00000000 ;
			15'h0000690A : data <= 8'b00000000 ;
			15'h0000690B : data <= 8'b00000000 ;
			15'h0000690C : data <= 8'b00000000 ;
			15'h0000690D : data <= 8'b00000000 ;
			15'h0000690E : data <= 8'b00000000 ;
			15'h0000690F : data <= 8'b00000000 ;
			15'h00006910 : data <= 8'b00000000 ;
			15'h00006911 : data <= 8'b00000000 ;
			15'h00006912 : data <= 8'b00000000 ;
			15'h00006913 : data <= 8'b00000000 ;
			15'h00006914 : data <= 8'b00000000 ;
			15'h00006915 : data <= 8'b00000000 ;
			15'h00006916 : data <= 8'b00000000 ;
			15'h00006917 : data <= 8'b00000000 ;
			15'h00006918 : data <= 8'b00000000 ;
			15'h00006919 : data <= 8'b00000000 ;
			15'h0000691A : data <= 8'b00000000 ;
			15'h0000691B : data <= 8'b00000000 ;
			15'h0000691C : data <= 8'b00000000 ;
			15'h0000691D : data <= 8'b00000000 ;
			15'h0000691E : data <= 8'b00000000 ;
			15'h0000691F : data <= 8'b00000000 ;
			15'h00006920 : data <= 8'b00000000 ;
			15'h00006921 : data <= 8'b00000000 ;
			15'h00006922 : data <= 8'b00000000 ;
			15'h00006923 : data <= 8'b00000000 ;
			15'h00006924 : data <= 8'b00000000 ;
			15'h00006925 : data <= 8'b00000000 ;
			15'h00006926 : data <= 8'b00000000 ;
			15'h00006927 : data <= 8'b00000000 ;
			15'h00006928 : data <= 8'b00000000 ;
			15'h00006929 : data <= 8'b00000000 ;
			15'h0000692A : data <= 8'b00000000 ;
			15'h0000692B : data <= 8'b00000000 ;
			15'h0000692C : data <= 8'b00000000 ;
			15'h0000692D : data <= 8'b00000000 ;
			15'h0000692E : data <= 8'b00000000 ;
			15'h0000692F : data <= 8'b00000000 ;
			15'h00006930 : data <= 8'b00000000 ;
			15'h00006931 : data <= 8'b00000000 ;
			15'h00006932 : data <= 8'b00000000 ;
			15'h00006933 : data <= 8'b00000000 ;
			15'h00006934 : data <= 8'b00000000 ;
			15'h00006935 : data <= 8'b00000000 ;
			15'h00006936 : data <= 8'b00000000 ;
			15'h00006937 : data <= 8'b00000000 ;
			15'h00006938 : data <= 8'b00000000 ;
			15'h00006939 : data <= 8'b00000000 ;
			15'h0000693A : data <= 8'b00000000 ;
			15'h0000693B : data <= 8'b00000000 ;
			15'h0000693C : data <= 8'b00000000 ;
			15'h0000693D : data <= 8'b00000000 ;
			15'h0000693E : data <= 8'b00000000 ;
			15'h0000693F : data <= 8'b00000000 ;
			15'h00006940 : data <= 8'b00000000 ;
			15'h00006941 : data <= 8'b00000000 ;
			15'h00006942 : data <= 8'b00000000 ;
			15'h00006943 : data <= 8'b00000000 ;
			15'h00006944 : data <= 8'b00000000 ;
			15'h00006945 : data <= 8'b00000000 ;
			15'h00006946 : data <= 8'b00000000 ;
			15'h00006947 : data <= 8'b00000000 ;
			15'h00006948 : data <= 8'b00000000 ;
			15'h00006949 : data <= 8'b00000000 ;
			15'h0000694A : data <= 8'b00000000 ;
			15'h0000694B : data <= 8'b00000000 ;
			15'h0000694C : data <= 8'b00000000 ;
			15'h0000694D : data <= 8'b00000000 ;
			15'h0000694E : data <= 8'b00000000 ;
			15'h0000694F : data <= 8'b00000000 ;
			15'h00006950 : data <= 8'b00000000 ;
			15'h00006951 : data <= 8'b00000000 ;
			15'h00006952 : data <= 8'b00000000 ;
			15'h00006953 : data <= 8'b00000000 ;
			15'h00006954 : data <= 8'b00000000 ;
			15'h00006955 : data <= 8'b00000000 ;
			15'h00006956 : data <= 8'b00000000 ;
			15'h00006957 : data <= 8'b00000000 ;
			15'h00006958 : data <= 8'b00000000 ;
			15'h00006959 : data <= 8'b00000000 ;
			15'h0000695A : data <= 8'b00000000 ;
			15'h0000695B : data <= 8'b00000000 ;
			15'h0000695C : data <= 8'b00000000 ;
			15'h0000695D : data <= 8'b00000000 ;
			15'h0000695E : data <= 8'b00000000 ;
			15'h0000695F : data <= 8'b00000000 ;
			15'h00006960 : data <= 8'b00000000 ;
			15'h00006961 : data <= 8'b00000000 ;
			15'h00006962 : data <= 8'b00000000 ;
			15'h00006963 : data <= 8'b00000000 ;
			15'h00006964 : data <= 8'b00000000 ;
			15'h00006965 : data <= 8'b00000000 ;
			15'h00006966 : data <= 8'b00000000 ;
			15'h00006967 : data <= 8'b00000000 ;
			15'h00006968 : data <= 8'b00000000 ;
			15'h00006969 : data <= 8'b00000000 ;
			15'h0000696A : data <= 8'b00000000 ;
			15'h0000696B : data <= 8'b00000000 ;
			15'h0000696C : data <= 8'b00000000 ;
			15'h0000696D : data <= 8'b00000000 ;
			15'h0000696E : data <= 8'b00000000 ;
			15'h0000696F : data <= 8'b00000000 ;
			15'h00006970 : data <= 8'b00000000 ;
			15'h00006971 : data <= 8'b00000000 ;
			15'h00006972 : data <= 8'b00000000 ;
			15'h00006973 : data <= 8'b00000000 ;
			15'h00006974 : data <= 8'b00000000 ;
			15'h00006975 : data <= 8'b00000000 ;
			15'h00006976 : data <= 8'b00000000 ;
			15'h00006977 : data <= 8'b00000000 ;
			15'h00006978 : data <= 8'b00000000 ;
			15'h00006979 : data <= 8'b00000000 ;
			15'h0000697A : data <= 8'b00000000 ;
			15'h0000697B : data <= 8'b00000000 ;
			15'h0000697C : data <= 8'b00000000 ;
			15'h0000697D : data <= 8'b00000000 ;
			15'h0000697E : data <= 8'b00000000 ;
			15'h0000697F : data <= 8'b00000000 ;
			15'h00006980 : data <= 8'b00000000 ;
			15'h00006981 : data <= 8'b00000000 ;
			15'h00006982 : data <= 8'b00000000 ;
			15'h00006983 : data <= 8'b00000000 ;
			15'h00006984 : data <= 8'b00000000 ;
			15'h00006985 : data <= 8'b00000000 ;
			15'h00006986 : data <= 8'b00000000 ;
			15'h00006987 : data <= 8'b00000000 ;
			15'h00006988 : data <= 8'b00000000 ;
			15'h00006989 : data <= 8'b00000000 ;
			15'h0000698A : data <= 8'b00000000 ;
			15'h0000698B : data <= 8'b00000000 ;
			15'h0000698C : data <= 8'b00000000 ;
			15'h0000698D : data <= 8'b00000000 ;
			15'h0000698E : data <= 8'b00000000 ;
			15'h0000698F : data <= 8'b00000000 ;
			15'h00006990 : data <= 8'b00000000 ;
			15'h00006991 : data <= 8'b00000000 ;
			15'h00006992 : data <= 8'b00000000 ;
			15'h00006993 : data <= 8'b00000000 ;
			15'h00006994 : data <= 8'b00000000 ;
			15'h00006995 : data <= 8'b00000000 ;
			15'h00006996 : data <= 8'b00000000 ;
			15'h00006997 : data <= 8'b00000000 ;
			15'h00006998 : data <= 8'b00000000 ;
			15'h00006999 : data <= 8'b00000000 ;
			15'h0000699A : data <= 8'b00000000 ;
			15'h0000699B : data <= 8'b00000000 ;
			15'h0000699C : data <= 8'b00000000 ;
			15'h0000699D : data <= 8'b00000000 ;
			15'h0000699E : data <= 8'b00000000 ;
			15'h0000699F : data <= 8'b00000000 ;
			15'h000069A0 : data <= 8'b00000000 ;
			15'h000069A1 : data <= 8'b00000000 ;
			15'h000069A2 : data <= 8'b00000000 ;
			15'h000069A3 : data <= 8'b00000000 ;
			15'h000069A4 : data <= 8'b00000000 ;
			15'h000069A5 : data <= 8'b00000000 ;
			15'h000069A6 : data <= 8'b00000000 ;
			15'h000069A7 : data <= 8'b00000000 ;
			15'h000069A8 : data <= 8'b00000000 ;
			15'h000069A9 : data <= 8'b00000000 ;
			15'h000069AA : data <= 8'b00000000 ;
			15'h000069AB : data <= 8'b00000000 ;
			15'h000069AC : data <= 8'b00000000 ;
			15'h000069AD : data <= 8'b00000000 ;
			15'h000069AE : data <= 8'b00000000 ;
			15'h000069AF : data <= 8'b00000000 ;
			15'h000069B0 : data <= 8'b00000000 ;
			15'h000069B1 : data <= 8'b00000000 ;
			15'h000069B2 : data <= 8'b00000000 ;
			15'h000069B3 : data <= 8'b00000000 ;
			15'h000069B4 : data <= 8'b00000000 ;
			15'h000069B5 : data <= 8'b00000000 ;
			15'h000069B6 : data <= 8'b00000000 ;
			15'h000069B7 : data <= 8'b00000000 ;
			15'h000069B8 : data <= 8'b00000000 ;
			15'h000069B9 : data <= 8'b00000000 ;
			15'h000069BA : data <= 8'b00000000 ;
			15'h000069BB : data <= 8'b00000000 ;
			15'h000069BC : data <= 8'b00000000 ;
			15'h000069BD : data <= 8'b00000000 ;
			15'h000069BE : data <= 8'b00000000 ;
			15'h000069BF : data <= 8'b00000000 ;
			15'h000069C0 : data <= 8'b00000000 ;
			15'h000069C1 : data <= 8'b00000000 ;
			15'h000069C2 : data <= 8'b00000000 ;
			15'h000069C3 : data <= 8'b00000000 ;
			15'h000069C4 : data <= 8'b00000000 ;
			15'h000069C5 : data <= 8'b00000000 ;
			15'h000069C6 : data <= 8'b00000000 ;
			15'h000069C7 : data <= 8'b00000000 ;
			15'h000069C8 : data <= 8'b00000000 ;
			15'h000069C9 : data <= 8'b00000000 ;
			15'h000069CA : data <= 8'b00000000 ;
			15'h000069CB : data <= 8'b00000000 ;
			15'h000069CC : data <= 8'b00000000 ;
			15'h000069CD : data <= 8'b00000000 ;
			15'h000069CE : data <= 8'b00000000 ;
			15'h000069CF : data <= 8'b00000000 ;
			15'h000069D0 : data <= 8'b00000000 ;
			15'h000069D1 : data <= 8'b00000000 ;
			15'h000069D2 : data <= 8'b00000000 ;
			15'h000069D3 : data <= 8'b00000000 ;
			15'h000069D4 : data <= 8'b00000000 ;
			15'h000069D5 : data <= 8'b00000000 ;
			15'h000069D6 : data <= 8'b00000000 ;
			15'h000069D7 : data <= 8'b00000000 ;
			15'h000069D8 : data <= 8'b00000000 ;
			15'h000069D9 : data <= 8'b00000000 ;
			15'h000069DA : data <= 8'b00000000 ;
			15'h000069DB : data <= 8'b00000000 ;
			15'h000069DC : data <= 8'b00000000 ;
			15'h000069DD : data <= 8'b00000000 ;
			15'h000069DE : data <= 8'b00000000 ;
			15'h000069DF : data <= 8'b00000000 ;
			15'h000069E0 : data <= 8'b00000000 ;
			15'h000069E1 : data <= 8'b00000000 ;
			15'h000069E2 : data <= 8'b00000000 ;
			15'h000069E3 : data <= 8'b00000000 ;
			15'h000069E4 : data <= 8'b00000000 ;
			15'h000069E5 : data <= 8'b00000000 ;
			15'h000069E6 : data <= 8'b00000000 ;
			15'h000069E7 : data <= 8'b00000000 ;
			15'h000069E8 : data <= 8'b00000000 ;
			15'h000069E9 : data <= 8'b00000000 ;
			15'h000069EA : data <= 8'b00000000 ;
			15'h000069EB : data <= 8'b00000000 ;
			15'h000069EC : data <= 8'b00000000 ;
			15'h000069ED : data <= 8'b00000000 ;
			15'h000069EE : data <= 8'b00000000 ;
			15'h000069EF : data <= 8'b00000000 ;
			15'h000069F0 : data <= 8'b00000000 ;
			15'h000069F1 : data <= 8'b00000000 ;
			15'h000069F2 : data <= 8'b00000000 ;
			15'h000069F3 : data <= 8'b00000000 ;
			15'h000069F4 : data <= 8'b00000000 ;
			15'h000069F5 : data <= 8'b00000000 ;
			15'h000069F6 : data <= 8'b00000000 ;
			15'h000069F7 : data <= 8'b00000000 ;
			15'h000069F8 : data <= 8'b00000000 ;
			15'h000069F9 : data <= 8'b00000000 ;
			15'h000069FA : data <= 8'b00000000 ;
			15'h000069FB : data <= 8'b00000000 ;
			15'h000069FC : data <= 8'b00000000 ;
			15'h000069FD : data <= 8'b00000000 ;
			15'h000069FE : data <= 8'b00000000 ;
			15'h000069FF : data <= 8'b00000000 ;
			15'h00006A00 : data <= 8'b00000000 ;
			15'h00006A01 : data <= 8'b00000000 ;
			15'h00006A02 : data <= 8'b00000000 ;
			15'h00006A03 : data <= 8'b00000000 ;
			15'h00006A04 : data <= 8'b00000000 ;
			15'h00006A05 : data <= 8'b00000000 ;
			15'h00006A06 : data <= 8'b00000000 ;
			15'h00006A07 : data <= 8'b00000000 ;
			15'h00006A08 : data <= 8'b00000000 ;
			15'h00006A09 : data <= 8'b00000000 ;
			15'h00006A0A : data <= 8'b00000000 ;
			15'h00006A0B : data <= 8'b00000000 ;
			15'h00006A0C : data <= 8'b00000000 ;
			15'h00006A0D : data <= 8'b00000000 ;
			15'h00006A0E : data <= 8'b00000000 ;
			15'h00006A0F : data <= 8'b00000000 ;
			15'h00006A10 : data <= 8'b00000000 ;
			15'h00006A11 : data <= 8'b00000000 ;
			15'h00006A12 : data <= 8'b00000000 ;
			15'h00006A13 : data <= 8'b00000000 ;
			15'h00006A14 : data <= 8'b00000000 ;
			15'h00006A15 : data <= 8'b00000000 ;
			15'h00006A16 : data <= 8'b00000000 ;
			15'h00006A17 : data <= 8'b00000000 ;
			15'h00006A18 : data <= 8'b00000000 ;
			15'h00006A19 : data <= 8'b00000000 ;
			15'h00006A1A : data <= 8'b00000000 ;
			15'h00006A1B : data <= 8'b00000000 ;
			15'h00006A1C : data <= 8'b00000000 ;
			15'h00006A1D : data <= 8'b00000000 ;
			15'h00006A1E : data <= 8'b00000000 ;
			15'h00006A1F : data <= 8'b00000000 ;
			15'h00006A20 : data <= 8'b00000000 ;
			15'h00006A21 : data <= 8'b00000000 ;
			15'h00006A22 : data <= 8'b00000000 ;
			15'h00006A23 : data <= 8'b00000000 ;
			15'h00006A24 : data <= 8'b00000000 ;
			15'h00006A25 : data <= 8'b00000000 ;
			15'h00006A26 : data <= 8'b00000000 ;
			15'h00006A27 : data <= 8'b00000000 ;
			15'h00006A28 : data <= 8'b00000000 ;
			15'h00006A29 : data <= 8'b00000000 ;
			15'h00006A2A : data <= 8'b00000000 ;
			15'h00006A2B : data <= 8'b00000000 ;
			15'h00006A2C : data <= 8'b00000000 ;
			15'h00006A2D : data <= 8'b00000000 ;
			15'h00006A2E : data <= 8'b00000000 ;
			15'h00006A2F : data <= 8'b00000000 ;
			15'h00006A30 : data <= 8'b00000000 ;
			15'h00006A31 : data <= 8'b00000000 ;
			15'h00006A32 : data <= 8'b00000000 ;
			15'h00006A33 : data <= 8'b00000000 ;
			15'h00006A34 : data <= 8'b00000000 ;
			15'h00006A35 : data <= 8'b00000000 ;
			15'h00006A36 : data <= 8'b00000000 ;
			15'h00006A37 : data <= 8'b00000000 ;
			15'h00006A38 : data <= 8'b00000000 ;
			15'h00006A39 : data <= 8'b00000000 ;
			15'h00006A3A : data <= 8'b00000000 ;
			15'h00006A3B : data <= 8'b00000000 ;
			15'h00006A3C : data <= 8'b00000000 ;
			15'h00006A3D : data <= 8'b00000000 ;
			15'h00006A3E : data <= 8'b00000000 ;
			15'h00006A3F : data <= 8'b00000000 ;
			15'h00006A40 : data <= 8'b00000000 ;
			15'h00006A41 : data <= 8'b00000000 ;
			15'h00006A42 : data <= 8'b00000000 ;
			15'h00006A43 : data <= 8'b00000000 ;
			15'h00006A44 : data <= 8'b00000000 ;
			15'h00006A45 : data <= 8'b00000000 ;
			15'h00006A46 : data <= 8'b00000000 ;
			15'h00006A47 : data <= 8'b00000000 ;
			15'h00006A48 : data <= 8'b00000000 ;
			15'h00006A49 : data <= 8'b00000000 ;
			15'h00006A4A : data <= 8'b00000000 ;
			15'h00006A4B : data <= 8'b00000000 ;
			15'h00006A4C : data <= 8'b00000000 ;
			15'h00006A4D : data <= 8'b00000000 ;
			15'h00006A4E : data <= 8'b00000000 ;
			15'h00006A4F : data <= 8'b00000000 ;
			15'h00006A50 : data <= 8'b00000000 ;
			15'h00006A51 : data <= 8'b00000000 ;
			15'h00006A52 : data <= 8'b00000000 ;
			15'h00006A53 : data <= 8'b00000000 ;
			15'h00006A54 : data <= 8'b00000000 ;
			15'h00006A55 : data <= 8'b00000000 ;
			15'h00006A56 : data <= 8'b00000000 ;
			15'h00006A57 : data <= 8'b00000000 ;
			15'h00006A58 : data <= 8'b00000000 ;
			15'h00006A59 : data <= 8'b00000000 ;
			15'h00006A5A : data <= 8'b00000000 ;
			15'h00006A5B : data <= 8'b00000000 ;
			15'h00006A5C : data <= 8'b00000000 ;
			15'h00006A5D : data <= 8'b00000000 ;
			15'h00006A5E : data <= 8'b00000000 ;
			15'h00006A5F : data <= 8'b00000000 ;
			15'h00006A60 : data <= 8'b00000000 ;
			15'h00006A61 : data <= 8'b00000000 ;
			15'h00006A62 : data <= 8'b00000000 ;
			15'h00006A63 : data <= 8'b00000000 ;
			15'h00006A64 : data <= 8'b00000000 ;
			15'h00006A65 : data <= 8'b00000000 ;
			15'h00006A66 : data <= 8'b00000000 ;
			15'h00006A67 : data <= 8'b00000000 ;
			15'h00006A68 : data <= 8'b00000000 ;
			15'h00006A69 : data <= 8'b00000000 ;
			15'h00006A6A : data <= 8'b00000000 ;
			15'h00006A6B : data <= 8'b00000000 ;
			15'h00006A6C : data <= 8'b00000000 ;
			15'h00006A6D : data <= 8'b00000000 ;
			15'h00006A6E : data <= 8'b00000000 ;
			15'h00006A6F : data <= 8'b00000000 ;
			15'h00006A70 : data <= 8'b00000000 ;
			15'h00006A71 : data <= 8'b00000000 ;
			15'h00006A72 : data <= 8'b00000000 ;
			15'h00006A73 : data <= 8'b00000000 ;
			15'h00006A74 : data <= 8'b00000000 ;
			15'h00006A75 : data <= 8'b00000000 ;
			15'h00006A76 : data <= 8'b00000000 ;
			15'h00006A77 : data <= 8'b00000000 ;
			15'h00006A78 : data <= 8'b00000000 ;
			15'h00006A79 : data <= 8'b00000000 ;
			15'h00006A7A : data <= 8'b00000000 ;
			15'h00006A7B : data <= 8'b00000000 ;
			15'h00006A7C : data <= 8'b00000000 ;
			15'h00006A7D : data <= 8'b00000000 ;
			15'h00006A7E : data <= 8'b00000000 ;
			15'h00006A7F : data <= 8'b00000000 ;
			15'h00006A80 : data <= 8'b00000000 ;
			15'h00006A81 : data <= 8'b00000000 ;
			15'h00006A82 : data <= 8'b00000000 ;
			15'h00006A83 : data <= 8'b00000000 ;
			15'h00006A84 : data <= 8'b00000000 ;
			15'h00006A85 : data <= 8'b00000000 ;
			15'h00006A86 : data <= 8'b00000000 ;
			15'h00006A87 : data <= 8'b00000000 ;
			15'h00006A88 : data <= 8'b00000000 ;
			15'h00006A89 : data <= 8'b00000000 ;
			15'h00006A8A : data <= 8'b00000000 ;
			15'h00006A8B : data <= 8'b00000000 ;
			15'h00006A8C : data <= 8'b00000000 ;
			15'h00006A8D : data <= 8'b00000000 ;
			15'h00006A8E : data <= 8'b00000000 ;
			15'h00006A8F : data <= 8'b00000000 ;
			15'h00006A90 : data <= 8'b00000000 ;
			15'h00006A91 : data <= 8'b00000000 ;
			15'h00006A92 : data <= 8'b00000000 ;
			15'h00006A93 : data <= 8'b00000000 ;
			15'h00006A94 : data <= 8'b00000000 ;
			15'h00006A95 : data <= 8'b00000000 ;
			15'h00006A96 : data <= 8'b00000000 ;
			15'h00006A97 : data <= 8'b00000000 ;
			15'h00006A98 : data <= 8'b00000000 ;
			15'h00006A99 : data <= 8'b00000000 ;
			15'h00006A9A : data <= 8'b00000000 ;
			15'h00006A9B : data <= 8'b00000000 ;
			15'h00006A9C : data <= 8'b00000000 ;
			15'h00006A9D : data <= 8'b00000000 ;
			15'h00006A9E : data <= 8'b00000000 ;
			15'h00006A9F : data <= 8'b00000000 ;
			15'h00006AA0 : data <= 8'b00000000 ;
			15'h00006AA1 : data <= 8'b00000000 ;
			15'h00006AA2 : data <= 8'b00000000 ;
			15'h00006AA3 : data <= 8'b00000000 ;
			15'h00006AA4 : data <= 8'b00000000 ;
			15'h00006AA5 : data <= 8'b00000000 ;
			15'h00006AA6 : data <= 8'b00000000 ;
			15'h00006AA7 : data <= 8'b00000000 ;
			15'h00006AA8 : data <= 8'b00000000 ;
			15'h00006AA9 : data <= 8'b00000000 ;
			15'h00006AAA : data <= 8'b00000000 ;
			15'h00006AAB : data <= 8'b00000000 ;
			15'h00006AAC : data <= 8'b00000000 ;
			15'h00006AAD : data <= 8'b00000000 ;
			15'h00006AAE : data <= 8'b00000000 ;
			15'h00006AAF : data <= 8'b00000000 ;
			15'h00006AB0 : data <= 8'b00000000 ;
			15'h00006AB1 : data <= 8'b00000000 ;
			15'h00006AB2 : data <= 8'b00000000 ;
			15'h00006AB3 : data <= 8'b00000000 ;
			15'h00006AB4 : data <= 8'b00000000 ;
			15'h00006AB5 : data <= 8'b00000000 ;
			15'h00006AB6 : data <= 8'b00000000 ;
			15'h00006AB7 : data <= 8'b00000000 ;
			15'h00006AB8 : data <= 8'b00000000 ;
			15'h00006AB9 : data <= 8'b00000000 ;
			15'h00006ABA : data <= 8'b00000000 ;
			15'h00006ABB : data <= 8'b00000000 ;
			15'h00006ABC : data <= 8'b00000000 ;
			15'h00006ABD : data <= 8'b00000000 ;
			15'h00006ABE : data <= 8'b00000000 ;
			15'h00006ABF : data <= 8'b00000000 ;
			15'h00006AC0 : data <= 8'b00000000 ;
			15'h00006AC1 : data <= 8'b00000000 ;
			15'h00006AC2 : data <= 8'b00000000 ;
			15'h00006AC3 : data <= 8'b00000000 ;
			15'h00006AC4 : data <= 8'b00000000 ;
			15'h00006AC5 : data <= 8'b00000000 ;
			15'h00006AC6 : data <= 8'b00000000 ;
			15'h00006AC7 : data <= 8'b00000000 ;
			15'h00006AC8 : data <= 8'b00000000 ;
			15'h00006AC9 : data <= 8'b00000000 ;
			15'h00006ACA : data <= 8'b00000000 ;
			15'h00006ACB : data <= 8'b00000000 ;
			15'h00006ACC : data <= 8'b00000000 ;
			15'h00006ACD : data <= 8'b00000000 ;
			15'h00006ACE : data <= 8'b00000000 ;
			15'h00006ACF : data <= 8'b00000000 ;
			15'h00006AD0 : data <= 8'b00000000 ;
			15'h00006AD1 : data <= 8'b00000000 ;
			15'h00006AD2 : data <= 8'b00000000 ;
			15'h00006AD3 : data <= 8'b00000000 ;
			15'h00006AD4 : data <= 8'b00000000 ;
			15'h00006AD5 : data <= 8'b00000000 ;
			15'h00006AD6 : data <= 8'b00000000 ;
			15'h00006AD7 : data <= 8'b00000000 ;
			15'h00006AD8 : data <= 8'b00000000 ;
			15'h00006AD9 : data <= 8'b00000000 ;
			15'h00006ADA : data <= 8'b00000000 ;
			15'h00006ADB : data <= 8'b00000000 ;
			15'h00006ADC : data <= 8'b00000000 ;
			15'h00006ADD : data <= 8'b00000000 ;
			15'h00006ADE : data <= 8'b00000000 ;
			15'h00006ADF : data <= 8'b00000000 ;
			15'h00006AE0 : data <= 8'b00000000 ;
			15'h00006AE1 : data <= 8'b00000000 ;
			15'h00006AE2 : data <= 8'b00000000 ;
			15'h00006AE3 : data <= 8'b00000000 ;
			15'h00006AE4 : data <= 8'b00000000 ;
			15'h00006AE5 : data <= 8'b00000000 ;
			15'h00006AE6 : data <= 8'b00000000 ;
			15'h00006AE7 : data <= 8'b00000000 ;
			15'h00006AE8 : data <= 8'b00000000 ;
			15'h00006AE9 : data <= 8'b00000000 ;
			15'h00006AEA : data <= 8'b00000000 ;
			15'h00006AEB : data <= 8'b00000000 ;
			15'h00006AEC : data <= 8'b00000000 ;
			15'h00006AED : data <= 8'b00000000 ;
			15'h00006AEE : data <= 8'b00000000 ;
			15'h00006AEF : data <= 8'b00000000 ;
			15'h00006AF0 : data <= 8'b00000000 ;
			15'h00006AF1 : data <= 8'b00000000 ;
			15'h00006AF2 : data <= 8'b00000000 ;
			15'h00006AF3 : data <= 8'b00000000 ;
			15'h00006AF4 : data <= 8'b00000000 ;
			15'h00006AF5 : data <= 8'b00000000 ;
			15'h00006AF6 : data <= 8'b00000000 ;
			15'h00006AF7 : data <= 8'b00000000 ;
			15'h00006AF8 : data <= 8'b00000000 ;
			15'h00006AF9 : data <= 8'b00000000 ;
			15'h00006AFA : data <= 8'b00000000 ;
			15'h00006AFB : data <= 8'b00000000 ;
			15'h00006AFC : data <= 8'b00000000 ;
			15'h00006AFD : data <= 8'b00000000 ;
			15'h00006AFE : data <= 8'b00000000 ;
			15'h00006AFF : data <= 8'b00000000 ;
			15'h00006B00 : data <= 8'b00000000 ;
			15'h00006B01 : data <= 8'b00000000 ;
			15'h00006B02 : data <= 8'b00000000 ;
			15'h00006B03 : data <= 8'b00000000 ;
			15'h00006B04 : data <= 8'b00000000 ;
			15'h00006B05 : data <= 8'b00000000 ;
			15'h00006B06 : data <= 8'b00000000 ;
			15'h00006B07 : data <= 8'b00000000 ;
			15'h00006B08 : data <= 8'b00000000 ;
			15'h00006B09 : data <= 8'b00000000 ;
			15'h00006B0A : data <= 8'b00000000 ;
			15'h00006B0B : data <= 8'b00000000 ;
			15'h00006B0C : data <= 8'b00000000 ;
			15'h00006B0D : data <= 8'b00000000 ;
			15'h00006B0E : data <= 8'b00000000 ;
			15'h00006B0F : data <= 8'b00000000 ;
			15'h00006B10 : data <= 8'b00000000 ;
			15'h00006B11 : data <= 8'b00000000 ;
			15'h00006B12 : data <= 8'b00000000 ;
			15'h00006B13 : data <= 8'b00000000 ;
			15'h00006B14 : data <= 8'b00000000 ;
			15'h00006B15 : data <= 8'b00000000 ;
			15'h00006B16 : data <= 8'b00000000 ;
			15'h00006B17 : data <= 8'b00000000 ;
			15'h00006B18 : data <= 8'b00000000 ;
			15'h00006B19 : data <= 8'b00000000 ;
			15'h00006B1A : data <= 8'b00000000 ;
			15'h00006B1B : data <= 8'b00000000 ;
			15'h00006B1C : data <= 8'b00000000 ;
			15'h00006B1D : data <= 8'b00000000 ;
			15'h00006B1E : data <= 8'b00000000 ;
			15'h00006B1F : data <= 8'b00000000 ;
			15'h00006B20 : data <= 8'b00000000 ;
			15'h00006B21 : data <= 8'b00000000 ;
			15'h00006B22 : data <= 8'b00000000 ;
			15'h00006B23 : data <= 8'b00000000 ;
			15'h00006B24 : data <= 8'b00000000 ;
			15'h00006B25 : data <= 8'b00000000 ;
			15'h00006B26 : data <= 8'b00000000 ;
			15'h00006B27 : data <= 8'b00000000 ;
			15'h00006B28 : data <= 8'b00000000 ;
			15'h00006B29 : data <= 8'b00000000 ;
			15'h00006B2A : data <= 8'b00000000 ;
			15'h00006B2B : data <= 8'b00000000 ;
			15'h00006B2C : data <= 8'b00000000 ;
			15'h00006B2D : data <= 8'b00000000 ;
			15'h00006B2E : data <= 8'b00000000 ;
			15'h00006B2F : data <= 8'b00000000 ;
			15'h00006B30 : data <= 8'b00000000 ;
			15'h00006B31 : data <= 8'b00000000 ;
			15'h00006B32 : data <= 8'b00000000 ;
			15'h00006B33 : data <= 8'b00000000 ;
			15'h00006B34 : data <= 8'b00000000 ;
			15'h00006B35 : data <= 8'b00000000 ;
			15'h00006B36 : data <= 8'b00000000 ;
			15'h00006B37 : data <= 8'b00000000 ;
			15'h00006B38 : data <= 8'b00000000 ;
			15'h00006B39 : data <= 8'b00000000 ;
			15'h00006B3A : data <= 8'b00000000 ;
			15'h00006B3B : data <= 8'b00000000 ;
			15'h00006B3C : data <= 8'b00000000 ;
			15'h00006B3D : data <= 8'b00000000 ;
			15'h00006B3E : data <= 8'b00000000 ;
			15'h00006B3F : data <= 8'b00000000 ;
			15'h00006B40 : data <= 8'b00000000 ;
			15'h00006B41 : data <= 8'b00000000 ;
			15'h00006B42 : data <= 8'b00000000 ;
			15'h00006B43 : data <= 8'b00000000 ;
			15'h00006B44 : data <= 8'b00000000 ;
			15'h00006B45 : data <= 8'b00000000 ;
			15'h00006B46 : data <= 8'b00000000 ;
			15'h00006B47 : data <= 8'b00000000 ;
			15'h00006B48 : data <= 8'b00000000 ;
			15'h00006B49 : data <= 8'b00000000 ;
			15'h00006B4A : data <= 8'b00000000 ;
			15'h00006B4B : data <= 8'b00000000 ;
			15'h00006B4C : data <= 8'b00000000 ;
			15'h00006B4D : data <= 8'b00000000 ;
			15'h00006B4E : data <= 8'b00000000 ;
			15'h00006B4F : data <= 8'b00000000 ;
			15'h00006B50 : data <= 8'b00000000 ;
			15'h00006B51 : data <= 8'b00000000 ;
			15'h00006B52 : data <= 8'b00000000 ;
			15'h00006B53 : data <= 8'b00000000 ;
			15'h00006B54 : data <= 8'b00000000 ;
			15'h00006B55 : data <= 8'b00000000 ;
			15'h00006B56 : data <= 8'b00000000 ;
			15'h00006B57 : data <= 8'b00000000 ;
			15'h00006B58 : data <= 8'b00000000 ;
			15'h00006B59 : data <= 8'b00000000 ;
			15'h00006B5A : data <= 8'b00000000 ;
			15'h00006B5B : data <= 8'b00000000 ;
			15'h00006B5C : data <= 8'b00000000 ;
			15'h00006B5D : data <= 8'b00000000 ;
			15'h00006B5E : data <= 8'b00000000 ;
			15'h00006B5F : data <= 8'b00000000 ;
			15'h00006B60 : data <= 8'b00000000 ;
			15'h00006B61 : data <= 8'b00000000 ;
			15'h00006B62 : data <= 8'b00000000 ;
			15'h00006B63 : data <= 8'b00000000 ;
			15'h00006B64 : data <= 8'b00000000 ;
			15'h00006B65 : data <= 8'b00000000 ;
			15'h00006B66 : data <= 8'b00000000 ;
			15'h00006B67 : data <= 8'b00000000 ;
			15'h00006B68 : data <= 8'b00000000 ;
			15'h00006B69 : data <= 8'b00000000 ;
			15'h00006B6A : data <= 8'b00000000 ;
			15'h00006B6B : data <= 8'b00000000 ;
			15'h00006B6C : data <= 8'b00000000 ;
			15'h00006B6D : data <= 8'b00000000 ;
			15'h00006B6E : data <= 8'b00000000 ;
			15'h00006B6F : data <= 8'b00000000 ;
			15'h00006B70 : data <= 8'b00000000 ;
			15'h00006B71 : data <= 8'b00000000 ;
			15'h00006B72 : data <= 8'b00000000 ;
			15'h00006B73 : data <= 8'b00000000 ;
			15'h00006B74 : data <= 8'b00000000 ;
			15'h00006B75 : data <= 8'b00000000 ;
			15'h00006B76 : data <= 8'b00000000 ;
			15'h00006B77 : data <= 8'b00000000 ;
			15'h00006B78 : data <= 8'b00000000 ;
			15'h00006B79 : data <= 8'b00000000 ;
			15'h00006B7A : data <= 8'b00000000 ;
			15'h00006B7B : data <= 8'b00000000 ;
			15'h00006B7C : data <= 8'b00000000 ;
			15'h00006B7D : data <= 8'b00000000 ;
			15'h00006B7E : data <= 8'b00000000 ;
			15'h00006B7F : data <= 8'b00000000 ;
			15'h00006B80 : data <= 8'b00000000 ;
			15'h00006B81 : data <= 8'b00000000 ;
			15'h00006B82 : data <= 8'b00000000 ;
			15'h00006B83 : data <= 8'b00000000 ;
			15'h00006B84 : data <= 8'b00000000 ;
			15'h00006B85 : data <= 8'b00000000 ;
			15'h00006B86 : data <= 8'b00000000 ;
			15'h00006B87 : data <= 8'b00000000 ;
			15'h00006B88 : data <= 8'b00000000 ;
			15'h00006B89 : data <= 8'b00000000 ;
			15'h00006B8A : data <= 8'b00000000 ;
			15'h00006B8B : data <= 8'b00000000 ;
			15'h00006B8C : data <= 8'b00000000 ;
			15'h00006B8D : data <= 8'b00000000 ;
			15'h00006B8E : data <= 8'b00000000 ;
			15'h00006B8F : data <= 8'b00000000 ;
			15'h00006B90 : data <= 8'b00000000 ;
			15'h00006B91 : data <= 8'b00000000 ;
			15'h00006B92 : data <= 8'b00000000 ;
			15'h00006B93 : data <= 8'b00000000 ;
			15'h00006B94 : data <= 8'b00000000 ;
			15'h00006B95 : data <= 8'b00000000 ;
			15'h00006B96 : data <= 8'b00000000 ;
			15'h00006B97 : data <= 8'b00000000 ;
			15'h00006B98 : data <= 8'b00000000 ;
			15'h00006B99 : data <= 8'b00000000 ;
			15'h00006B9A : data <= 8'b00000000 ;
			15'h00006B9B : data <= 8'b00000000 ;
			15'h00006B9C : data <= 8'b00000000 ;
			15'h00006B9D : data <= 8'b00000000 ;
			15'h00006B9E : data <= 8'b00000000 ;
			15'h00006B9F : data <= 8'b00000000 ;
			15'h00006BA0 : data <= 8'b00000000 ;
			15'h00006BA1 : data <= 8'b00000000 ;
			15'h00006BA2 : data <= 8'b00000000 ;
			15'h00006BA3 : data <= 8'b00000000 ;
			15'h00006BA4 : data <= 8'b00000000 ;
			15'h00006BA5 : data <= 8'b00000000 ;
			15'h00006BA6 : data <= 8'b00000000 ;
			15'h00006BA7 : data <= 8'b00000000 ;
			15'h00006BA8 : data <= 8'b00000000 ;
			15'h00006BA9 : data <= 8'b00000000 ;
			15'h00006BAA : data <= 8'b00000000 ;
			15'h00006BAB : data <= 8'b00000000 ;
			15'h00006BAC : data <= 8'b00000000 ;
			15'h00006BAD : data <= 8'b00000000 ;
			15'h00006BAE : data <= 8'b00000000 ;
			15'h00006BAF : data <= 8'b00000000 ;
			15'h00006BB0 : data <= 8'b00000000 ;
			15'h00006BB1 : data <= 8'b00000000 ;
			15'h00006BB2 : data <= 8'b00000000 ;
			15'h00006BB3 : data <= 8'b00000000 ;
			15'h00006BB4 : data <= 8'b00000000 ;
			15'h00006BB5 : data <= 8'b00000000 ;
			15'h00006BB6 : data <= 8'b00000000 ;
			15'h00006BB7 : data <= 8'b00000000 ;
			15'h00006BB8 : data <= 8'b00000000 ;
			15'h00006BB9 : data <= 8'b00000000 ;
			15'h00006BBA : data <= 8'b00000000 ;
			15'h00006BBB : data <= 8'b00000000 ;
			15'h00006BBC : data <= 8'b00000000 ;
			15'h00006BBD : data <= 8'b00000000 ;
			15'h00006BBE : data <= 8'b00000000 ;
			15'h00006BBF : data <= 8'b00000000 ;
			15'h00006BC0 : data <= 8'b00000000 ;
			15'h00006BC1 : data <= 8'b00000000 ;
			15'h00006BC2 : data <= 8'b00000000 ;
			15'h00006BC3 : data <= 8'b00000000 ;
			15'h00006BC4 : data <= 8'b00000000 ;
			15'h00006BC5 : data <= 8'b00000000 ;
			15'h00006BC6 : data <= 8'b00000000 ;
			15'h00006BC7 : data <= 8'b00000000 ;
			15'h00006BC8 : data <= 8'b00000000 ;
			15'h00006BC9 : data <= 8'b00000000 ;
			15'h00006BCA : data <= 8'b00000000 ;
			15'h00006BCB : data <= 8'b00000000 ;
			15'h00006BCC : data <= 8'b00000000 ;
			15'h00006BCD : data <= 8'b00000000 ;
			15'h00006BCE : data <= 8'b00000000 ;
			15'h00006BCF : data <= 8'b00000000 ;
			15'h00006BD0 : data <= 8'b00000000 ;
			15'h00006BD1 : data <= 8'b00000000 ;
			15'h00006BD2 : data <= 8'b00000000 ;
			15'h00006BD3 : data <= 8'b00000000 ;
			15'h00006BD4 : data <= 8'b00000000 ;
			15'h00006BD5 : data <= 8'b00000000 ;
			15'h00006BD6 : data <= 8'b00000000 ;
			15'h00006BD7 : data <= 8'b00000000 ;
			15'h00006BD8 : data <= 8'b00000000 ;
			15'h00006BD9 : data <= 8'b00000000 ;
			15'h00006BDA : data <= 8'b00000000 ;
			15'h00006BDB : data <= 8'b00000000 ;
			15'h00006BDC : data <= 8'b00000000 ;
			15'h00006BDD : data <= 8'b00000000 ;
			15'h00006BDE : data <= 8'b00000000 ;
			15'h00006BDF : data <= 8'b00000000 ;
			15'h00006BE0 : data <= 8'b00000000 ;
			15'h00006BE1 : data <= 8'b00000000 ;
			15'h00006BE2 : data <= 8'b00000000 ;
			15'h00006BE3 : data <= 8'b00000000 ;
			15'h00006BE4 : data <= 8'b00000000 ;
			15'h00006BE5 : data <= 8'b00000000 ;
			15'h00006BE6 : data <= 8'b00000000 ;
			15'h00006BE7 : data <= 8'b00000000 ;
			15'h00006BE8 : data <= 8'b00000000 ;
			15'h00006BE9 : data <= 8'b00000000 ;
			15'h00006BEA : data <= 8'b00000000 ;
			15'h00006BEB : data <= 8'b00000000 ;
			15'h00006BEC : data <= 8'b00000000 ;
			15'h00006BED : data <= 8'b00000000 ;
			15'h00006BEE : data <= 8'b00000000 ;
			15'h00006BEF : data <= 8'b00000000 ;
			15'h00006BF0 : data <= 8'b00000000 ;
			15'h00006BF1 : data <= 8'b00000000 ;
			15'h00006BF2 : data <= 8'b00000000 ;
			15'h00006BF3 : data <= 8'b00000000 ;
			15'h00006BF4 : data <= 8'b00000000 ;
			15'h00006BF5 : data <= 8'b00000000 ;
			15'h00006BF6 : data <= 8'b00000000 ;
			15'h00006BF7 : data <= 8'b00000000 ;
			15'h00006BF8 : data <= 8'b00000000 ;
			15'h00006BF9 : data <= 8'b00000000 ;
			15'h00006BFA : data <= 8'b00000000 ;
			15'h00006BFB : data <= 8'b00000000 ;
			15'h00006BFC : data <= 8'b00000000 ;
			15'h00006BFD : data <= 8'b00000000 ;
			15'h00006BFE : data <= 8'b00000000 ;
			15'h00006BFF : data <= 8'b00000000 ;
			15'h00006C00 : data <= 8'b00000000 ;
			15'h00006C01 : data <= 8'b00000000 ;
			15'h00006C02 : data <= 8'b00000000 ;
			15'h00006C03 : data <= 8'b00000000 ;
			15'h00006C04 : data <= 8'b00000000 ;
			15'h00006C05 : data <= 8'b00000000 ;
			15'h00006C06 : data <= 8'b00000000 ;
			15'h00006C07 : data <= 8'b00000000 ;
			15'h00006C08 : data <= 8'b00000000 ;
			15'h00006C09 : data <= 8'b00000000 ;
			15'h00006C0A : data <= 8'b00000000 ;
			15'h00006C0B : data <= 8'b00000000 ;
			15'h00006C0C : data <= 8'b00000000 ;
			15'h00006C0D : data <= 8'b00000000 ;
			15'h00006C0E : data <= 8'b00000000 ;
			15'h00006C0F : data <= 8'b00000000 ;
			15'h00006C10 : data <= 8'b00000000 ;
			15'h00006C11 : data <= 8'b00000000 ;
			15'h00006C12 : data <= 8'b00000000 ;
			15'h00006C13 : data <= 8'b00000000 ;
			15'h00006C14 : data <= 8'b00000000 ;
			15'h00006C15 : data <= 8'b00000000 ;
			15'h00006C16 : data <= 8'b00000000 ;
			15'h00006C17 : data <= 8'b00000000 ;
			15'h00006C18 : data <= 8'b00000000 ;
			15'h00006C19 : data <= 8'b00000000 ;
			15'h00006C1A : data <= 8'b00000000 ;
			15'h00006C1B : data <= 8'b00000000 ;
			15'h00006C1C : data <= 8'b00000000 ;
			15'h00006C1D : data <= 8'b00000000 ;
			15'h00006C1E : data <= 8'b00000000 ;
			15'h00006C1F : data <= 8'b00000000 ;
			15'h00006C20 : data <= 8'b00000000 ;
			15'h00006C21 : data <= 8'b00000000 ;
			15'h00006C22 : data <= 8'b00000000 ;
			15'h00006C23 : data <= 8'b00000000 ;
			15'h00006C24 : data <= 8'b00000000 ;
			15'h00006C25 : data <= 8'b00000000 ;
			15'h00006C26 : data <= 8'b00000000 ;
			15'h00006C27 : data <= 8'b00000000 ;
			15'h00006C28 : data <= 8'b00000000 ;
			15'h00006C29 : data <= 8'b00000000 ;
			15'h00006C2A : data <= 8'b00000000 ;
			15'h00006C2B : data <= 8'b00000000 ;
			15'h00006C2C : data <= 8'b00000000 ;
			15'h00006C2D : data <= 8'b00000000 ;
			15'h00006C2E : data <= 8'b00000000 ;
			15'h00006C2F : data <= 8'b00000000 ;
			15'h00006C30 : data <= 8'b00000000 ;
			15'h00006C31 : data <= 8'b00000000 ;
			15'h00006C32 : data <= 8'b00000000 ;
			15'h00006C33 : data <= 8'b00000000 ;
			15'h00006C34 : data <= 8'b00000000 ;
			15'h00006C35 : data <= 8'b00000000 ;
			15'h00006C36 : data <= 8'b00000000 ;
			15'h00006C37 : data <= 8'b00000000 ;
			15'h00006C38 : data <= 8'b00000000 ;
			15'h00006C39 : data <= 8'b00000000 ;
			15'h00006C3A : data <= 8'b00000000 ;
			15'h00006C3B : data <= 8'b00000000 ;
			15'h00006C3C : data <= 8'b00000000 ;
			15'h00006C3D : data <= 8'b00000000 ;
			15'h00006C3E : data <= 8'b00000000 ;
			15'h00006C3F : data <= 8'b00000000 ;
			15'h00006C40 : data <= 8'b00000000 ;
			15'h00006C41 : data <= 8'b00000000 ;
			15'h00006C42 : data <= 8'b00000000 ;
			15'h00006C43 : data <= 8'b00000000 ;
			15'h00006C44 : data <= 8'b00000000 ;
			15'h00006C45 : data <= 8'b00000000 ;
			15'h00006C46 : data <= 8'b00000000 ;
			15'h00006C47 : data <= 8'b00000000 ;
			15'h00006C48 : data <= 8'b00000000 ;
			15'h00006C49 : data <= 8'b00000000 ;
			15'h00006C4A : data <= 8'b00000000 ;
			15'h00006C4B : data <= 8'b00000000 ;
			15'h00006C4C : data <= 8'b00000000 ;
			15'h00006C4D : data <= 8'b00000000 ;
			15'h00006C4E : data <= 8'b00000000 ;
			15'h00006C4F : data <= 8'b00000000 ;
			15'h00006C50 : data <= 8'b00000000 ;
			15'h00006C51 : data <= 8'b00000000 ;
			15'h00006C52 : data <= 8'b00000000 ;
			15'h00006C53 : data <= 8'b00000000 ;
			15'h00006C54 : data <= 8'b00000000 ;
			15'h00006C55 : data <= 8'b00000000 ;
			15'h00006C56 : data <= 8'b00000000 ;
			15'h00006C57 : data <= 8'b00000000 ;
			15'h00006C58 : data <= 8'b00000000 ;
			15'h00006C59 : data <= 8'b00000000 ;
			15'h00006C5A : data <= 8'b00000000 ;
			15'h00006C5B : data <= 8'b00000000 ;
			15'h00006C5C : data <= 8'b00000000 ;
			15'h00006C5D : data <= 8'b00000000 ;
			15'h00006C5E : data <= 8'b00000000 ;
			15'h00006C5F : data <= 8'b00000000 ;
			15'h00006C60 : data <= 8'b00000000 ;
			15'h00006C61 : data <= 8'b00000000 ;
			15'h00006C62 : data <= 8'b00000000 ;
			15'h00006C63 : data <= 8'b00000000 ;
			15'h00006C64 : data <= 8'b00000000 ;
			15'h00006C65 : data <= 8'b00000000 ;
			15'h00006C66 : data <= 8'b00000000 ;
			15'h00006C67 : data <= 8'b00000000 ;
			15'h00006C68 : data <= 8'b00000000 ;
			15'h00006C69 : data <= 8'b00000000 ;
			15'h00006C6A : data <= 8'b00000000 ;
			15'h00006C6B : data <= 8'b00000000 ;
			15'h00006C6C : data <= 8'b00000000 ;
			15'h00006C6D : data <= 8'b00000000 ;
			15'h00006C6E : data <= 8'b00000000 ;
			15'h00006C6F : data <= 8'b00000000 ;
			15'h00006C70 : data <= 8'b00000000 ;
			15'h00006C71 : data <= 8'b00000000 ;
			15'h00006C72 : data <= 8'b00000000 ;
			15'h00006C73 : data <= 8'b00000000 ;
			15'h00006C74 : data <= 8'b00000000 ;
			15'h00006C75 : data <= 8'b00000000 ;
			15'h00006C76 : data <= 8'b00000000 ;
			15'h00006C77 : data <= 8'b00000000 ;
			15'h00006C78 : data <= 8'b00000000 ;
			15'h00006C79 : data <= 8'b00000000 ;
			15'h00006C7A : data <= 8'b00000000 ;
			15'h00006C7B : data <= 8'b00000000 ;
			15'h00006C7C : data <= 8'b00000000 ;
			15'h00006C7D : data <= 8'b00000000 ;
			15'h00006C7E : data <= 8'b00000000 ;
			15'h00006C7F : data <= 8'b00000000 ;
			15'h00006C80 : data <= 8'b00000000 ;
			15'h00006C81 : data <= 8'b00000000 ;
			15'h00006C82 : data <= 8'b00000000 ;
			15'h00006C83 : data <= 8'b00000000 ;
			15'h00006C84 : data <= 8'b00000000 ;
			15'h00006C85 : data <= 8'b00000000 ;
			15'h00006C86 : data <= 8'b00000000 ;
			15'h00006C87 : data <= 8'b00000000 ;
			15'h00006C88 : data <= 8'b00000000 ;
			15'h00006C89 : data <= 8'b00000000 ;
			15'h00006C8A : data <= 8'b00000000 ;
			15'h00006C8B : data <= 8'b00000000 ;
			15'h00006C8C : data <= 8'b00000000 ;
			15'h00006C8D : data <= 8'b00000000 ;
			15'h00006C8E : data <= 8'b00000000 ;
			15'h00006C8F : data <= 8'b00000000 ;
			15'h00006C90 : data <= 8'b00000000 ;
			15'h00006C91 : data <= 8'b00000000 ;
			15'h00006C92 : data <= 8'b00000000 ;
			15'h00006C93 : data <= 8'b00000000 ;
			15'h00006C94 : data <= 8'b00000000 ;
			15'h00006C95 : data <= 8'b00000000 ;
			15'h00006C96 : data <= 8'b00000000 ;
			15'h00006C97 : data <= 8'b00000000 ;
			15'h00006C98 : data <= 8'b00000000 ;
			15'h00006C99 : data <= 8'b00000000 ;
			15'h00006C9A : data <= 8'b00000000 ;
			15'h00006C9B : data <= 8'b00000000 ;
			15'h00006C9C : data <= 8'b00000000 ;
			15'h00006C9D : data <= 8'b00000000 ;
			15'h00006C9E : data <= 8'b00000000 ;
			15'h00006C9F : data <= 8'b00000000 ;
			15'h00006CA0 : data <= 8'b00000000 ;
			15'h00006CA1 : data <= 8'b00000000 ;
			15'h00006CA2 : data <= 8'b00000000 ;
			15'h00006CA3 : data <= 8'b00000000 ;
			15'h00006CA4 : data <= 8'b00000000 ;
			15'h00006CA5 : data <= 8'b00000000 ;
			15'h00006CA6 : data <= 8'b00000000 ;
			15'h00006CA7 : data <= 8'b00000000 ;
			15'h00006CA8 : data <= 8'b00000000 ;
			15'h00006CA9 : data <= 8'b00000000 ;
			15'h00006CAA : data <= 8'b00000000 ;
			15'h00006CAB : data <= 8'b00000000 ;
			15'h00006CAC : data <= 8'b00000000 ;
			15'h00006CAD : data <= 8'b00000000 ;
			15'h00006CAE : data <= 8'b00000000 ;
			15'h00006CAF : data <= 8'b00000000 ;
			15'h00006CB0 : data <= 8'b00000000 ;
			15'h00006CB1 : data <= 8'b00000000 ;
			15'h00006CB2 : data <= 8'b00000000 ;
			15'h00006CB3 : data <= 8'b00000000 ;
			15'h00006CB4 : data <= 8'b00000000 ;
			15'h00006CB5 : data <= 8'b00000000 ;
			15'h00006CB6 : data <= 8'b00000000 ;
			15'h00006CB7 : data <= 8'b00000000 ;
			15'h00006CB8 : data <= 8'b00000000 ;
			15'h00006CB9 : data <= 8'b00000000 ;
			15'h00006CBA : data <= 8'b00000000 ;
			15'h00006CBB : data <= 8'b00000000 ;
			15'h00006CBC : data <= 8'b00000000 ;
			15'h00006CBD : data <= 8'b00000000 ;
			15'h00006CBE : data <= 8'b00000000 ;
			15'h00006CBF : data <= 8'b00000000 ;
			15'h00006CC0 : data <= 8'b00000000 ;
			15'h00006CC1 : data <= 8'b00000000 ;
			15'h00006CC2 : data <= 8'b00000000 ;
			15'h00006CC3 : data <= 8'b00000000 ;
			15'h00006CC4 : data <= 8'b00000000 ;
			15'h00006CC5 : data <= 8'b00000000 ;
			15'h00006CC6 : data <= 8'b00000000 ;
			15'h00006CC7 : data <= 8'b00000000 ;
			15'h00006CC8 : data <= 8'b00000000 ;
			15'h00006CC9 : data <= 8'b00000000 ;
			15'h00006CCA : data <= 8'b00000000 ;
			15'h00006CCB : data <= 8'b00000000 ;
			15'h00006CCC : data <= 8'b00000000 ;
			15'h00006CCD : data <= 8'b00000000 ;
			15'h00006CCE : data <= 8'b00000000 ;
			15'h00006CCF : data <= 8'b00000000 ;
			15'h00006CD0 : data <= 8'b00000000 ;
			15'h00006CD1 : data <= 8'b00000000 ;
			15'h00006CD2 : data <= 8'b00000000 ;
			15'h00006CD3 : data <= 8'b00000000 ;
			15'h00006CD4 : data <= 8'b00000000 ;
			15'h00006CD5 : data <= 8'b00000000 ;
			15'h00006CD6 : data <= 8'b00000000 ;
			15'h00006CD7 : data <= 8'b00000000 ;
			15'h00006CD8 : data <= 8'b00000000 ;
			15'h00006CD9 : data <= 8'b00000000 ;
			15'h00006CDA : data <= 8'b00000000 ;
			15'h00006CDB : data <= 8'b00000000 ;
			15'h00006CDC : data <= 8'b00000000 ;
			15'h00006CDD : data <= 8'b00000000 ;
			15'h00006CDE : data <= 8'b00000000 ;
			15'h00006CDF : data <= 8'b00000000 ;
			15'h00006CE0 : data <= 8'b00000000 ;
			15'h00006CE1 : data <= 8'b00000000 ;
			15'h00006CE2 : data <= 8'b00000000 ;
			15'h00006CE3 : data <= 8'b00000000 ;
			15'h00006CE4 : data <= 8'b00000000 ;
			15'h00006CE5 : data <= 8'b00000000 ;
			15'h00006CE6 : data <= 8'b00000000 ;
			15'h00006CE7 : data <= 8'b00000000 ;
			15'h00006CE8 : data <= 8'b00000000 ;
			15'h00006CE9 : data <= 8'b00000000 ;
			15'h00006CEA : data <= 8'b00000000 ;
			15'h00006CEB : data <= 8'b00000000 ;
			15'h00006CEC : data <= 8'b00000000 ;
			15'h00006CED : data <= 8'b00000000 ;
			15'h00006CEE : data <= 8'b00000000 ;
			15'h00006CEF : data <= 8'b00000000 ;
			15'h00006CF0 : data <= 8'b00000000 ;
			15'h00006CF1 : data <= 8'b00000000 ;
			15'h00006CF2 : data <= 8'b00000000 ;
			15'h00006CF3 : data <= 8'b00000000 ;
			15'h00006CF4 : data <= 8'b00000000 ;
			15'h00006CF5 : data <= 8'b00000000 ;
			15'h00006CF6 : data <= 8'b00000000 ;
			15'h00006CF7 : data <= 8'b00000000 ;
			15'h00006CF8 : data <= 8'b00000000 ;
			15'h00006CF9 : data <= 8'b00000000 ;
			15'h00006CFA : data <= 8'b00000000 ;
			15'h00006CFB : data <= 8'b00000000 ;
			15'h00006CFC : data <= 8'b00000000 ;
			15'h00006CFD : data <= 8'b00000000 ;
			15'h00006CFE : data <= 8'b00000000 ;
			15'h00006CFF : data <= 8'b00000000 ;
			15'h00006D00 : data <= 8'b00000000 ;
			15'h00006D01 : data <= 8'b00000000 ;
			15'h00006D02 : data <= 8'b00000000 ;
			15'h00006D03 : data <= 8'b00000000 ;
			15'h00006D04 : data <= 8'b00000000 ;
			15'h00006D05 : data <= 8'b00000000 ;
			15'h00006D06 : data <= 8'b00000000 ;
			15'h00006D07 : data <= 8'b00000000 ;
			15'h00006D08 : data <= 8'b00000000 ;
			15'h00006D09 : data <= 8'b00000000 ;
			15'h00006D0A : data <= 8'b00000000 ;
			15'h00006D0B : data <= 8'b00000000 ;
			15'h00006D0C : data <= 8'b00000000 ;
			15'h00006D0D : data <= 8'b00000000 ;
			15'h00006D0E : data <= 8'b00000000 ;
			15'h00006D0F : data <= 8'b00000000 ;
			15'h00006D10 : data <= 8'b00000000 ;
			15'h00006D11 : data <= 8'b00000000 ;
			15'h00006D12 : data <= 8'b00000000 ;
			15'h00006D13 : data <= 8'b00000000 ;
			15'h00006D14 : data <= 8'b00000000 ;
			15'h00006D15 : data <= 8'b00000000 ;
			15'h00006D16 : data <= 8'b00000000 ;
			15'h00006D17 : data <= 8'b00000000 ;
			15'h00006D18 : data <= 8'b00000000 ;
			15'h00006D19 : data <= 8'b00000000 ;
			15'h00006D1A : data <= 8'b00000000 ;
			15'h00006D1B : data <= 8'b00000000 ;
			15'h00006D1C : data <= 8'b00000000 ;
			15'h00006D1D : data <= 8'b00000000 ;
			15'h00006D1E : data <= 8'b00000000 ;
			15'h00006D1F : data <= 8'b00000000 ;
			15'h00006D20 : data <= 8'b00000000 ;
			15'h00006D21 : data <= 8'b00000000 ;
			15'h00006D22 : data <= 8'b00000000 ;
			15'h00006D23 : data <= 8'b00000000 ;
			15'h00006D24 : data <= 8'b00000000 ;
			15'h00006D25 : data <= 8'b00000000 ;
			15'h00006D26 : data <= 8'b00000000 ;
			15'h00006D27 : data <= 8'b00000000 ;
			15'h00006D28 : data <= 8'b00000000 ;
			15'h00006D29 : data <= 8'b00000000 ;
			15'h00006D2A : data <= 8'b00000000 ;
			15'h00006D2B : data <= 8'b00000000 ;
			15'h00006D2C : data <= 8'b00000000 ;
			15'h00006D2D : data <= 8'b00000000 ;
			15'h00006D2E : data <= 8'b00000000 ;
			15'h00006D2F : data <= 8'b00000000 ;
			15'h00006D30 : data <= 8'b00000000 ;
			15'h00006D31 : data <= 8'b00000000 ;
			15'h00006D32 : data <= 8'b00000000 ;
			15'h00006D33 : data <= 8'b00000000 ;
			15'h00006D34 : data <= 8'b00000000 ;
			15'h00006D35 : data <= 8'b00000000 ;
			15'h00006D36 : data <= 8'b00000000 ;
			15'h00006D37 : data <= 8'b00000000 ;
			15'h00006D38 : data <= 8'b00000000 ;
			15'h00006D39 : data <= 8'b00000000 ;
			15'h00006D3A : data <= 8'b00000000 ;
			15'h00006D3B : data <= 8'b00000000 ;
			15'h00006D3C : data <= 8'b00000000 ;
			15'h00006D3D : data <= 8'b00000000 ;
			15'h00006D3E : data <= 8'b00000000 ;
			15'h00006D3F : data <= 8'b00000000 ;
			15'h00006D40 : data <= 8'b00000000 ;
			15'h00006D41 : data <= 8'b00000000 ;
			15'h00006D42 : data <= 8'b00000000 ;
			15'h00006D43 : data <= 8'b00000000 ;
			15'h00006D44 : data <= 8'b00000000 ;
			15'h00006D45 : data <= 8'b00000000 ;
			15'h00006D46 : data <= 8'b00000000 ;
			15'h00006D47 : data <= 8'b00000000 ;
			15'h00006D48 : data <= 8'b00000000 ;
			15'h00006D49 : data <= 8'b00000000 ;
			15'h00006D4A : data <= 8'b00000000 ;
			15'h00006D4B : data <= 8'b00000000 ;
			15'h00006D4C : data <= 8'b00000000 ;
			15'h00006D4D : data <= 8'b00000000 ;
			15'h00006D4E : data <= 8'b00000000 ;
			15'h00006D4F : data <= 8'b00000000 ;
			15'h00006D50 : data <= 8'b00000000 ;
			15'h00006D51 : data <= 8'b00000000 ;
			15'h00006D52 : data <= 8'b00000000 ;
			15'h00006D53 : data <= 8'b00000000 ;
			15'h00006D54 : data <= 8'b00000000 ;
			15'h00006D55 : data <= 8'b00000000 ;
			15'h00006D56 : data <= 8'b00000000 ;
			15'h00006D57 : data <= 8'b00000000 ;
			15'h00006D58 : data <= 8'b00000000 ;
			15'h00006D59 : data <= 8'b00000000 ;
			15'h00006D5A : data <= 8'b00000000 ;
			15'h00006D5B : data <= 8'b00000000 ;
			15'h00006D5C : data <= 8'b00000000 ;
			15'h00006D5D : data <= 8'b00000000 ;
			15'h00006D5E : data <= 8'b00000000 ;
			15'h00006D5F : data <= 8'b00000000 ;
			15'h00006D60 : data <= 8'b00000000 ;
			15'h00006D61 : data <= 8'b00000000 ;
			15'h00006D62 : data <= 8'b00000000 ;
			15'h00006D63 : data <= 8'b00000000 ;
			15'h00006D64 : data <= 8'b00000000 ;
			15'h00006D65 : data <= 8'b00000000 ;
			15'h00006D66 : data <= 8'b00000000 ;
			15'h00006D67 : data <= 8'b00000000 ;
			15'h00006D68 : data <= 8'b00000000 ;
			15'h00006D69 : data <= 8'b00000000 ;
			15'h00006D6A : data <= 8'b00000000 ;
			15'h00006D6B : data <= 8'b00000000 ;
			15'h00006D6C : data <= 8'b00000000 ;
			15'h00006D6D : data <= 8'b00000000 ;
			15'h00006D6E : data <= 8'b00000000 ;
			15'h00006D6F : data <= 8'b00000000 ;
			15'h00006D70 : data <= 8'b00000000 ;
			15'h00006D71 : data <= 8'b00000000 ;
			15'h00006D72 : data <= 8'b00000000 ;
			15'h00006D73 : data <= 8'b00000000 ;
			15'h00006D74 : data <= 8'b00000000 ;
			15'h00006D75 : data <= 8'b00000000 ;
			15'h00006D76 : data <= 8'b00000000 ;
			15'h00006D77 : data <= 8'b00000000 ;
			15'h00006D78 : data <= 8'b00000000 ;
			15'h00006D79 : data <= 8'b00000000 ;
			15'h00006D7A : data <= 8'b00000000 ;
			15'h00006D7B : data <= 8'b00000000 ;
			15'h00006D7C : data <= 8'b00000000 ;
			15'h00006D7D : data <= 8'b00000000 ;
			15'h00006D7E : data <= 8'b00000000 ;
			15'h00006D7F : data <= 8'b00000000 ;
			15'h00006D80 : data <= 8'b00000000 ;
			15'h00006D81 : data <= 8'b00000000 ;
			15'h00006D82 : data <= 8'b00000000 ;
			15'h00006D83 : data <= 8'b00000000 ;
			15'h00006D84 : data <= 8'b00000000 ;
			15'h00006D85 : data <= 8'b00000000 ;
			15'h00006D86 : data <= 8'b00000000 ;
			15'h00006D87 : data <= 8'b00000000 ;
			15'h00006D88 : data <= 8'b00000000 ;
			15'h00006D89 : data <= 8'b00000000 ;
			15'h00006D8A : data <= 8'b00000000 ;
			15'h00006D8B : data <= 8'b00000000 ;
			15'h00006D8C : data <= 8'b00000000 ;
			15'h00006D8D : data <= 8'b00000000 ;
			15'h00006D8E : data <= 8'b00000000 ;
			15'h00006D8F : data <= 8'b00000000 ;
			15'h00006D90 : data <= 8'b00000000 ;
			15'h00006D91 : data <= 8'b00000000 ;
			15'h00006D92 : data <= 8'b00000000 ;
			15'h00006D93 : data <= 8'b00000000 ;
			15'h00006D94 : data <= 8'b00000000 ;
			15'h00006D95 : data <= 8'b00000000 ;
			15'h00006D96 : data <= 8'b00000000 ;
			15'h00006D97 : data <= 8'b00000000 ;
			15'h00006D98 : data <= 8'b00000000 ;
			15'h00006D99 : data <= 8'b00000000 ;
			15'h00006D9A : data <= 8'b00000000 ;
			15'h00006D9B : data <= 8'b00000000 ;
			15'h00006D9C : data <= 8'b00000000 ;
			15'h00006D9D : data <= 8'b00000000 ;
			15'h00006D9E : data <= 8'b00000000 ;
			15'h00006D9F : data <= 8'b00000000 ;
			15'h00006DA0 : data <= 8'b00000000 ;
			15'h00006DA1 : data <= 8'b00000000 ;
			15'h00006DA2 : data <= 8'b00000000 ;
			15'h00006DA3 : data <= 8'b00000000 ;
			15'h00006DA4 : data <= 8'b00000000 ;
			15'h00006DA5 : data <= 8'b00000000 ;
			15'h00006DA6 : data <= 8'b00000000 ;
			15'h00006DA7 : data <= 8'b00000000 ;
			15'h00006DA8 : data <= 8'b00000000 ;
			15'h00006DA9 : data <= 8'b00000000 ;
			15'h00006DAA : data <= 8'b00000000 ;
			15'h00006DAB : data <= 8'b00000000 ;
			15'h00006DAC : data <= 8'b00000000 ;
			15'h00006DAD : data <= 8'b00000000 ;
			15'h00006DAE : data <= 8'b00000000 ;
			15'h00006DAF : data <= 8'b00000000 ;
			15'h00006DB0 : data <= 8'b00000000 ;
			15'h00006DB1 : data <= 8'b00000000 ;
			15'h00006DB2 : data <= 8'b00000000 ;
			15'h00006DB3 : data <= 8'b00000000 ;
			15'h00006DB4 : data <= 8'b00000000 ;
			15'h00006DB5 : data <= 8'b00000000 ;
			15'h00006DB6 : data <= 8'b00000000 ;
			15'h00006DB7 : data <= 8'b00000000 ;
			15'h00006DB8 : data <= 8'b00000000 ;
			15'h00006DB9 : data <= 8'b00000000 ;
			15'h00006DBA : data <= 8'b00000000 ;
			15'h00006DBB : data <= 8'b00000000 ;
			15'h00006DBC : data <= 8'b00000000 ;
			15'h00006DBD : data <= 8'b00000000 ;
			15'h00006DBE : data <= 8'b00000000 ;
			15'h00006DBF : data <= 8'b00000000 ;
			15'h00006DC0 : data <= 8'b00000000 ;
			15'h00006DC1 : data <= 8'b00000000 ;
			15'h00006DC2 : data <= 8'b00000000 ;
			15'h00006DC3 : data <= 8'b00000000 ;
			15'h00006DC4 : data <= 8'b00000000 ;
			15'h00006DC5 : data <= 8'b00000000 ;
			15'h00006DC6 : data <= 8'b00000000 ;
			15'h00006DC7 : data <= 8'b00000000 ;
			15'h00006DC8 : data <= 8'b00000000 ;
			15'h00006DC9 : data <= 8'b00000000 ;
			15'h00006DCA : data <= 8'b00000000 ;
			15'h00006DCB : data <= 8'b00000000 ;
			15'h00006DCC : data <= 8'b00000000 ;
			15'h00006DCD : data <= 8'b00000000 ;
			15'h00006DCE : data <= 8'b00000000 ;
			15'h00006DCF : data <= 8'b00000000 ;
			15'h00006DD0 : data <= 8'b00000000 ;
			15'h00006DD1 : data <= 8'b00000000 ;
			15'h00006DD2 : data <= 8'b00000000 ;
			15'h00006DD3 : data <= 8'b00000000 ;
			15'h00006DD4 : data <= 8'b00000000 ;
			15'h00006DD5 : data <= 8'b00000000 ;
			15'h00006DD6 : data <= 8'b00000000 ;
			15'h00006DD7 : data <= 8'b00000000 ;
			15'h00006DD8 : data <= 8'b00000000 ;
			15'h00006DD9 : data <= 8'b00000000 ;
			15'h00006DDA : data <= 8'b00000000 ;
			15'h00006DDB : data <= 8'b00000000 ;
			15'h00006DDC : data <= 8'b00000000 ;
			15'h00006DDD : data <= 8'b00000000 ;
			15'h00006DDE : data <= 8'b00000000 ;
			15'h00006DDF : data <= 8'b00000000 ;
			15'h00006DE0 : data <= 8'b00000000 ;
			15'h00006DE1 : data <= 8'b00000000 ;
			15'h00006DE2 : data <= 8'b00000000 ;
			15'h00006DE3 : data <= 8'b00000000 ;
			15'h00006DE4 : data <= 8'b00000000 ;
			15'h00006DE5 : data <= 8'b00000000 ;
			15'h00006DE6 : data <= 8'b00000000 ;
			15'h00006DE7 : data <= 8'b00000000 ;
			15'h00006DE8 : data <= 8'b00000000 ;
			15'h00006DE9 : data <= 8'b00000000 ;
			15'h00006DEA : data <= 8'b00000000 ;
			15'h00006DEB : data <= 8'b00000000 ;
			15'h00006DEC : data <= 8'b00000000 ;
			15'h00006DED : data <= 8'b00000000 ;
			15'h00006DEE : data <= 8'b00000000 ;
			15'h00006DEF : data <= 8'b00000000 ;
			15'h00006DF0 : data <= 8'b00000000 ;
			15'h00006DF1 : data <= 8'b00000000 ;
			15'h00006DF2 : data <= 8'b00000000 ;
			15'h00006DF3 : data <= 8'b00000000 ;
			15'h00006DF4 : data <= 8'b00000000 ;
			15'h00006DF5 : data <= 8'b00000000 ;
			15'h00006DF6 : data <= 8'b00000000 ;
			15'h00006DF7 : data <= 8'b00000000 ;
			15'h00006DF8 : data <= 8'b00000000 ;
			15'h00006DF9 : data <= 8'b00000000 ;
			15'h00006DFA : data <= 8'b00000000 ;
			15'h00006DFB : data <= 8'b00000000 ;
			15'h00006DFC : data <= 8'b00000000 ;
			15'h00006DFD : data <= 8'b00000000 ;
			15'h00006DFE : data <= 8'b00000000 ;
			15'h00006DFF : data <= 8'b00000000 ;
			15'h00006E00 : data <= 8'b00000000 ;
			15'h00006E01 : data <= 8'b00000000 ;
			15'h00006E02 : data <= 8'b00000000 ;
			15'h00006E03 : data <= 8'b00000000 ;
			15'h00006E04 : data <= 8'b00000000 ;
			15'h00006E05 : data <= 8'b00000000 ;
			15'h00006E06 : data <= 8'b00000000 ;
			15'h00006E07 : data <= 8'b00000000 ;
			15'h00006E08 : data <= 8'b00000000 ;
			15'h00006E09 : data <= 8'b00000000 ;
			15'h00006E0A : data <= 8'b00000000 ;
			15'h00006E0B : data <= 8'b00000000 ;
			15'h00006E0C : data <= 8'b00000000 ;
			15'h00006E0D : data <= 8'b00000000 ;
			15'h00006E0E : data <= 8'b00000000 ;
			15'h00006E0F : data <= 8'b00000000 ;
			15'h00006E10 : data <= 8'b00000000 ;
			15'h00006E11 : data <= 8'b00000000 ;
			15'h00006E12 : data <= 8'b00000000 ;
			15'h00006E13 : data <= 8'b00000000 ;
			15'h00006E14 : data <= 8'b00000000 ;
			15'h00006E15 : data <= 8'b00000000 ;
			15'h00006E16 : data <= 8'b00000000 ;
			15'h00006E17 : data <= 8'b00000000 ;
			15'h00006E18 : data <= 8'b00000000 ;
			15'h00006E19 : data <= 8'b00000000 ;
			15'h00006E1A : data <= 8'b00000000 ;
			15'h00006E1B : data <= 8'b00000000 ;
			15'h00006E1C : data <= 8'b00000000 ;
			15'h00006E1D : data <= 8'b00000000 ;
			15'h00006E1E : data <= 8'b00000000 ;
			15'h00006E1F : data <= 8'b00000000 ;
			15'h00006E20 : data <= 8'b00000000 ;
			15'h00006E21 : data <= 8'b00000000 ;
			15'h00006E22 : data <= 8'b00000000 ;
			15'h00006E23 : data <= 8'b00000000 ;
			15'h00006E24 : data <= 8'b00000000 ;
			15'h00006E25 : data <= 8'b00000000 ;
			15'h00006E26 : data <= 8'b00000000 ;
			15'h00006E27 : data <= 8'b00000000 ;
			15'h00006E28 : data <= 8'b00000000 ;
			15'h00006E29 : data <= 8'b00000000 ;
			15'h00006E2A : data <= 8'b00000000 ;
			15'h00006E2B : data <= 8'b00000000 ;
			15'h00006E2C : data <= 8'b00000000 ;
			15'h00006E2D : data <= 8'b00000000 ;
			15'h00006E2E : data <= 8'b00000000 ;
			15'h00006E2F : data <= 8'b00000000 ;
			15'h00006E30 : data <= 8'b00000000 ;
			15'h00006E31 : data <= 8'b00000000 ;
			15'h00006E32 : data <= 8'b00000000 ;
			15'h00006E33 : data <= 8'b00000000 ;
			15'h00006E34 : data <= 8'b00000000 ;
			15'h00006E35 : data <= 8'b00000000 ;
			15'h00006E36 : data <= 8'b00000000 ;
			15'h00006E37 : data <= 8'b00000000 ;
			15'h00006E38 : data <= 8'b00000000 ;
			15'h00006E39 : data <= 8'b00000000 ;
			15'h00006E3A : data <= 8'b00000000 ;
			15'h00006E3B : data <= 8'b00000000 ;
			15'h00006E3C : data <= 8'b00000000 ;
			15'h00006E3D : data <= 8'b00000000 ;
			15'h00006E3E : data <= 8'b00000000 ;
			15'h00006E3F : data <= 8'b00000000 ;
			15'h00006E40 : data <= 8'b00000000 ;
			15'h00006E41 : data <= 8'b00000000 ;
			15'h00006E42 : data <= 8'b00000000 ;
			15'h00006E43 : data <= 8'b00000000 ;
			15'h00006E44 : data <= 8'b00000000 ;
			15'h00006E45 : data <= 8'b00000000 ;
			15'h00006E46 : data <= 8'b00000000 ;
			15'h00006E47 : data <= 8'b00000000 ;
			15'h00006E48 : data <= 8'b00000000 ;
			15'h00006E49 : data <= 8'b00000000 ;
			15'h00006E4A : data <= 8'b00000000 ;
			15'h00006E4B : data <= 8'b00000000 ;
			15'h00006E4C : data <= 8'b00000000 ;
			15'h00006E4D : data <= 8'b00000000 ;
			15'h00006E4E : data <= 8'b00000000 ;
			15'h00006E4F : data <= 8'b00000000 ;
			15'h00006E50 : data <= 8'b00000000 ;
			15'h00006E51 : data <= 8'b00000000 ;
			15'h00006E52 : data <= 8'b00000000 ;
			15'h00006E53 : data <= 8'b00000000 ;
			15'h00006E54 : data <= 8'b00000000 ;
			15'h00006E55 : data <= 8'b00000000 ;
			15'h00006E56 : data <= 8'b00000000 ;
			15'h00006E57 : data <= 8'b00000000 ;
			15'h00006E58 : data <= 8'b00000000 ;
			15'h00006E59 : data <= 8'b00000000 ;
			15'h00006E5A : data <= 8'b00000000 ;
			15'h00006E5B : data <= 8'b00000000 ;
			15'h00006E5C : data <= 8'b00000000 ;
			15'h00006E5D : data <= 8'b00000000 ;
			15'h00006E5E : data <= 8'b00000000 ;
			15'h00006E5F : data <= 8'b00000000 ;
			15'h00006E60 : data <= 8'b00000000 ;
			15'h00006E61 : data <= 8'b00000000 ;
			15'h00006E62 : data <= 8'b00000000 ;
			15'h00006E63 : data <= 8'b00000000 ;
			15'h00006E64 : data <= 8'b00000000 ;
			15'h00006E65 : data <= 8'b00000000 ;
			15'h00006E66 : data <= 8'b00000000 ;
			15'h00006E67 : data <= 8'b00000000 ;
			15'h00006E68 : data <= 8'b00000000 ;
			15'h00006E69 : data <= 8'b00000000 ;
			15'h00006E6A : data <= 8'b00000000 ;
			15'h00006E6B : data <= 8'b00000000 ;
			15'h00006E6C : data <= 8'b00000000 ;
			15'h00006E6D : data <= 8'b00000000 ;
			15'h00006E6E : data <= 8'b00000000 ;
			15'h00006E6F : data <= 8'b00000000 ;
			15'h00006E70 : data <= 8'b00000000 ;
			15'h00006E71 : data <= 8'b00000000 ;
			15'h00006E72 : data <= 8'b00000000 ;
			15'h00006E73 : data <= 8'b00000000 ;
			15'h00006E74 : data <= 8'b00000000 ;
			15'h00006E75 : data <= 8'b00000000 ;
			15'h00006E76 : data <= 8'b00000000 ;
			15'h00006E77 : data <= 8'b00000000 ;
			15'h00006E78 : data <= 8'b00000000 ;
			15'h00006E79 : data <= 8'b00000000 ;
			15'h00006E7A : data <= 8'b00000000 ;
			15'h00006E7B : data <= 8'b00000000 ;
			15'h00006E7C : data <= 8'b00000000 ;
			15'h00006E7D : data <= 8'b00000000 ;
			15'h00006E7E : data <= 8'b00000000 ;
			15'h00006E7F : data <= 8'b00000000 ;
			15'h00006E80 : data <= 8'b00000000 ;
			15'h00006E81 : data <= 8'b00000000 ;
			15'h00006E82 : data <= 8'b00000000 ;
			15'h00006E83 : data <= 8'b00000000 ;
			15'h00006E84 : data <= 8'b00000000 ;
			15'h00006E85 : data <= 8'b00000000 ;
			15'h00006E86 : data <= 8'b00000000 ;
			15'h00006E87 : data <= 8'b00000000 ;
			15'h00006E88 : data <= 8'b00000000 ;
			15'h00006E89 : data <= 8'b00000000 ;
			15'h00006E8A : data <= 8'b00000000 ;
			15'h00006E8B : data <= 8'b00000000 ;
			15'h00006E8C : data <= 8'b00000000 ;
			15'h00006E8D : data <= 8'b00000000 ;
			15'h00006E8E : data <= 8'b00000000 ;
			15'h00006E8F : data <= 8'b00000000 ;
			15'h00006E90 : data <= 8'b00000000 ;
			15'h00006E91 : data <= 8'b00000000 ;
			15'h00006E92 : data <= 8'b00000000 ;
			15'h00006E93 : data <= 8'b00000000 ;
			15'h00006E94 : data <= 8'b00000000 ;
			15'h00006E95 : data <= 8'b00000000 ;
			15'h00006E96 : data <= 8'b00000000 ;
			15'h00006E97 : data <= 8'b00000000 ;
			15'h00006E98 : data <= 8'b00000000 ;
			15'h00006E99 : data <= 8'b00000000 ;
			15'h00006E9A : data <= 8'b00000000 ;
			15'h00006E9B : data <= 8'b00000000 ;
			15'h00006E9C : data <= 8'b00000000 ;
			15'h00006E9D : data <= 8'b00000000 ;
			15'h00006E9E : data <= 8'b00000000 ;
			15'h00006E9F : data <= 8'b00000000 ;
			15'h00006EA0 : data <= 8'b00000000 ;
			15'h00006EA1 : data <= 8'b00000000 ;
			15'h00006EA2 : data <= 8'b00000000 ;
			15'h00006EA3 : data <= 8'b00000000 ;
			15'h00006EA4 : data <= 8'b00000000 ;
			15'h00006EA5 : data <= 8'b00000000 ;
			15'h00006EA6 : data <= 8'b00000000 ;
			15'h00006EA7 : data <= 8'b00000000 ;
			15'h00006EA8 : data <= 8'b00000000 ;
			15'h00006EA9 : data <= 8'b00000000 ;
			15'h00006EAA : data <= 8'b00000000 ;
			15'h00006EAB : data <= 8'b00000000 ;
			15'h00006EAC : data <= 8'b00000000 ;
			15'h00006EAD : data <= 8'b00000000 ;
			15'h00006EAE : data <= 8'b00000000 ;
			15'h00006EAF : data <= 8'b00000000 ;
			15'h00006EB0 : data <= 8'b00000000 ;
			15'h00006EB1 : data <= 8'b00000000 ;
			15'h00006EB2 : data <= 8'b00000000 ;
			15'h00006EB3 : data <= 8'b00000000 ;
			15'h00006EB4 : data <= 8'b00000000 ;
			15'h00006EB5 : data <= 8'b00000000 ;
			15'h00006EB6 : data <= 8'b00000000 ;
			15'h00006EB7 : data <= 8'b00000000 ;
			15'h00006EB8 : data <= 8'b00000000 ;
			15'h00006EB9 : data <= 8'b00000000 ;
			15'h00006EBA : data <= 8'b00000000 ;
			15'h00006EBB : data <= 8'b00000000 ;
			15'h00006EBC : data <= 8'b00000000 ;
			15'h00006EBD : data <= 8'b00000000 ;
			15'h00006EBE : data <= 8'b00000000 ;
			15'h00006EBF : data <= 8'b00000000 ;
			15'h00006EC0 : data <= 8'b00000000 ;
			15'h00006EC1 : data <= 8'b00000000 ;
			15'h00006EC2 : data <= 8'b00000000 ;
			15'h00006EC3 : data <= 8'b00000000 ;
			15'h00006EC4 : data <= 8'b00000000 ;
			15'h00006EC5 : data <= 8'b00000000 ;
			15'h00006EC6 : data <= 8'b00000000 ;
			15'h00006EC7 : data <= 8'b00000000 ;
			15'h00006EC8 : data <= 8'b00000000 ;
			15'h00006EC9 : data <= 8'b00000000 ;
			15'h00006ECA : data <= 8'b00000000 ;
			15'h00006ECB : data <= 8'b00000000 ;
			15'h00006ECC : data <= 8'b00000000 ;
			15'h00006ECD : data <= 8'b00000000 ;
			15'h00006ECE : data <= 8'b00000000 ;
			15'h00006ECF : data <= 8'b00000000 ;
			15'h00006ED0 : data <= 8'b00000000 ;
			15'h00006ED1 : data <= 8'b00000000 ;
			15'h00006ED2 : data <= 8'b00000000 ;
			15'h00006ED3 : data <= 8'b00000000 ;
			15'h00006ED4 : data <= 8'b00000000 ;
			15'h00006ED5 : data <= 8'b00000000 ;
			15'h00006ED6 : data <= 8'b00000000 ;
			15'h00006ED7 : data <= 8'b00000000 ;
			15'h00006ED8 : data <= 8'b00000000 ;
			15'h00006ED9 : data <= 8'b00000000 ;
			15'h00006EDA : data <= 8'b00000000 ;
			15'h00006EDB : data <= 8'b00000000 ;
			15'h00006EDC : data <= 8'b00000000 ;
			15'h00006EDD : data <= 8'b00000000 ;
			15'h00006EDE : data <= 8'b00000000 ;
			15'h00006EDF : data <= 8'b00000000 ;
			15'h00006EE0 : data <= 8'b00000000 ;
			15'h00006EE1 : data <= 8'b00000000 ;
			15'h00006EE2 : data <= 8'b00000000 ;
			15'h00006EE3 : data <= 8'b00000000 ;
			15'h00006EE4 : data <= 8'b00000000 ;
			15'h00006EE5 : data <= 8'b00000000 ;
			15'h00006EE6 : data <= 8'b00000000 ;
			15'h00006EE7 : data <= 8'b00000000 ;
			15'h00006EE8 : data <= 8'b00000000 ;
			15'h00006EE9 : data <= 8'b00000000 ;
			15'h00006EEA : data <= 8'b00000000 ;
			15'h00006EEB : data <= 8'b00000000 ;
			15'h00006EEC : data <= 8'b00000000 ;
			15'h00006EED : data <= 8'b00000000 ;
			15'h00006EEE : data <= 8'b00000000 ;
			15'h00006EEF : data <= 8'b00000000 ;
			15'h00006EF0 : data <= 8'b00000000 ;
			15'h00006EF1 : data <= 8'b00000000 ;
			15'h00006EF2 : data <= 8'b00000000 ;
			15'h00006EF3 : data <= 8'b00000000 ;
			15'h00006EF4 : data <= 8'b00000000 ;
			15'h00006EF5 : data <= 8'b00000000 ;
			15'h00006EF6 : data <= 8'b00000000 ;
			15'h00006EF7 : data <= 8'b00000000 ;
			15'h00006EF8 : data <= 8'b00000000 ;
			15'h00006EF9 : data <= 8'b00000000 ;
			15'h00006EFA : data <= 8'b00000000 ;
			15'h00006EFB : data <= 8'b00000000 ;
			15'h00006EFC : data <= 8'b00000000 ;
			15'h00006EFD : data <= 8'b00000000 ;
			15'h00006EFE : data <= 8'b00000000 ;
			15'h00006EFF : data <= 8'b00000000 ;
			15'h00006F00 : data <= 8'b00000000 ;
			15'h00006F01 : data <= 8'b00000000 ;
			15'h00006F02 : data <= 8'b00000000 ;
			15'h00006F03 : data <= 8'b00000000 ;
			15'h00006F04 : data <= 8'b00000000 ;
			15'h00006F05 : data <= 8'b00000000 ;
			15'h00006F06 : data <= 8'b00000000 ;
			15'h00006F07 : data <= 8'b00000000 ;
			15'h00006F08 : data <= 8'b00000000 ;
			15'h00006F09 : data <= 8'b00000000 ;
			15'h00006F0A : data <= 8'b00000000 ;
			15'h00006F0B : data <= 8'b00000000 ;
			15'h00006F0C : data <= 8'b00000000 ;
			15'h00006F0D : data <= 8'b00000000 ;
			15'h00006F0E : data <= 8'b00000000 ;
			15'h00006F0F : data <= 8'b00000000 ;
			15'h00006F10 : data <= 8'b00000000 ;
			15'h00006F11 : data <= 8'b00000000 ;
			15'h00006F12 : data <= 8'b00000000 ;
			15'h00006F13 : data <= 8'b00000000 ;
			15'h00006F14 : data <= 8'b00000000 ;
			15'h00006F15 : data <= 8'b00000000 ;
			15'h00006F16 : data <= 8'b00000000 ;
			15'h00006F17 : data <= 8'b00000000 ;
			15'h00006F18 : data <= 8'b00000000 ;
			15'h00006F19 : data <= 8'b00000000 ;
			15'h00006F1A : data <= 8'b00000000 ;
			15'h00006F1B : data <= 8'b00000000 ;
			15'h00006F1C : data <= 8'b00000000 ;
			15'h00006F1D : data <= 8'b00000000 ;
			15'h00006F1E : data <= 8'b00000000 ;
			15'h00006F1F : data <= 8'b00000000 ;
			15'h00006F20 : data <= 8'b00000000 ;
			15'h00006F21 : data <= 8'b00000000 ;
			15'h00006F22 : data <= 8'b00000000 ;
			15'h00006F23 : data <= 8'b00000000 ;
			15'h00006F24 : data <= 8'b00000000 ;
			15'h00006F25 : data <= 8'b00000000 ;
			15'h00006F26 : data <= 8'b00000000 ;
			15'h00006F27 : data <= 8'b00000000 ;
			15'h00006F28 : data <= 8'b00000000 ;
			15'h00006F29 : data <= 8'b00000000 ;
			15'h00006F2A : data <= 8'b00000000 ;
			15'h00006F2B : data <= 8'b00000000 ;
			15'h00006F2C : data <= 8'b00000000 ;
			15'h00006F2D : data <= 8'b00000000 ;
			15'h00006F2E : data <= 8'b00000000 ;
			15'h00006F2F : data <= 8'b00000000 ;
			15'h00006F30 : data <= 8'b00000000 ;
			15'h00006F31 : data <= 8'b00000000 ;
			15'h00006F32 : data <= 8'b00000000 ;
			15'h00006F33 : data <= 8'b00000000 ;
			15'h00006F34 : data <= 8'b00000000 ;
			15'h00006F35 : data <= 8'b00000000 ;
			15'h00006F36 : data <= 8'b00000000 ;
			15'h00006F37 : data <= 8'b00000000 ;
			15'h00006F38 : data <= 8'b00000000 ;
			15'h00006F39 : data <= 8'b00000000 ;
			15'h00006F3A : data <= 8'b00000000 ;
			15'h00006F3B : data <= 8'b00000000 ;
			15'h00006F3C : data <= 8'b00000000 ;
			15'h00006F3D : data <= 8'b00000000 ;
			15'h00006F3E : data <= 8'b00000000 ;
			15'h00006F3F : data <= 8'b00000000 ;
			15'h00006F40 : data <= 8'b00000000 ;
			15'h00006F41 : data <= 8'b00000000 ;
			15'h00006F42 : data <= 8'b00000000 ;
			15'h00006F43 : data <= 8'b00000000 ;
			15'h00006F44 : data <= 8'b00000000 ;
			15'h00006F45 : data <= 8'b00000000 ;
			15'h00006F46 : data <= 8'b00000000 ;
			15'h00006F47 : data <= 8'b00000000 ;
			15'h00006F48 : data <= 8'b00000000 ;
			15'h00006F49 : data <= 8'b00000000 ;
			15'h00006F4A : data <= 8'b00000000 ;
			15'h00006F4B : data <= 8'b00000000 ;
			15'h00006F4C : data <= 8'b00000000 ;
			15'h00006F4D : data <= 8'b00000000 ;
			15'h00006F4E : data <= 8'b00000000 ;
			15'h00006F4F : data <= 8'b00000000 ;
			15'h00006F50 : data <= 8'b00000000 ;
			15'h00006F51 : data <= 8'b00000000 ;
			15'h00006F52 : data <= 8'b00000000 ;
			15'h00006F53 : data <= 8'b00000000 ;
			15'h00006F54 : data <= 8'b00000000 ;
			15'h00006F55 : data <= 8'b00000000 ;
			15'h00006F56 : data <= 8'b00000000 ;
			15'h00006F57 : data <= 8'b00000000 ;
			15'h00006F58 : data <= 8'b00000000 ;
			15'h00006F59 : data <= 8'b00000000 ;
			15'h00006F5A : data <= 8'b00000000 ;
			15'h00006F5B : data <= 8'b00000000 ;
			15'h00006F5C : data <= 8'b00000000 ;
			15'h00006F5D : data <= 8'b00000000 ;
			15'h00006F5E : data <= 8'b00000000 ;
			15'h00006F5F : data <= 8'b00000000 ;
			15'h00006F60 : data <= 8'b00000000 ;
			15'h00006F61 : data <= 8'b00000000 ;
			15'h00006F62 : data <= 8'b00000000 ;
			15'h00006F63 : data <= 8'b00000000 ;
			15'h00006F64 : data <= 8'b00000000 ;
			15'h00006F65 : data <= 8'b00000000 ;
			15'h00006F66 : data <= 8'b00000000 ;
			15'h00006F67 : data <= 8'b00000000 ;
			15'h00006F68 : data <= 8'b00000000 ;
			15'h00006F69 : data <= 8'b00000000 ;
			15'h00006F6A : data <= 8'b00000000 ;
			15'h00006F6B : data <= 8'b00000000 ;
			15'h00006F6C : data <= 8'b00000000 ;
			15'h00006F6D : data <= 8'b00000000 ;
			15'h00006F6E : data <= 8'b00000000 ;
			15'h00006F6F : data <= 8'b00000000 ;
			15'h00006F70 : data <= 8'b00000000 ;
			15'h00006F71 : data <= 8'b00000000 ;
			15'h00006F72 : data <= 8'b00000000 ;
			15'h00006F73 : data <= 8'b00000000 ;
			15'h00006F74 : data <= 8'b00000000 ;
			15'h00006F75 : data <= 8'b00000000 ;
			15'h00006F76 : data <= 8'b00000000 ;
			15'h00006F77 : data <= 8'b00000000 ;
			15'h00006F78 : data <= 8'b00000000 ;
			15'h00006F79 : data <= 8'b00000000 ;
			15'h00006F7A : data <= 8'b00000000 ;
			15'h00006F7B : data <= 8'b00000000 ;
			15'h00006F7C : data <= 8'b00000000 ;
			15'h00006F7D : data <= 8'b00000000 ;
			15'h00006F7E : data <= 8'b00000000 ;
			15'h00006F7F : data <= 8'b00000000 ;
			15'h00006F80 : data <= 8'b00000000 ;
			15'h00006F81 : data <= 8'b00000000 ;
			15'h00006F82 : data <= 8'b00000000 ;
			15'h00006F83 : data <= 8'b00000000 ;
			15'h00006F84 : data <= 8'b00000000 ;
			15'h00006F85 : data <= 8'b00000000 ;
			15'h00006F86 : data <= 8'b00000000 ;
			15'h00006F87 : data <= 8'b00000000 ;
			15'h00006F88 : data <= 8'b00000000 ;
			15'h00006F89 : data <= 8'b00000000 ;
			15'h00006F8A : data <= 8'b00000000 ;
			15'h00006F8B : data <= 8'b00000000 ;
			15'h00006F8C : data <= 8'b00000000 ;
			15'h00006F8D : data <= 8'b00000000 ;
			15'h00006F8E : data <= 8'b00000000 ;
			15'h00006F8F : data <= 8'b00000000 ;
			15'h00006F90 : data <= 8'b00000000 ;
			15'h00006F91 : data <= 8'b00000000 ;
			15'h00006F92 : data <= 8'b00000000 ;
			15'h00006F93 : data <= 8'b00000000 ;
			15'h00006F94 : data <= 8'b00000000 ;
			15'h00006F95 : data <= 8'b00000000 ;
			15'h00006F96 : data <= 8'b00000000 ;
			15'h00006F97 : data <= 8'b00000000 ;
			15'h00006F98 : data <= 8'b00000000 ;
			15'h00006F99 : data <= 8'b00000000 ;
			15'h00006F9A : data <= 8'b00000000 ;
			15'h00006F9B : data <= 8'b00000000 ;
			15'h00006F9C : data <= 8'b00000000 ;
			15'h00006F9D : data <= 8'b00000000 ;
			15'h00006F9E : data <= 8'b00000000 ;
			15'h00006F9F : data <= 8'b00000000 ;
			15'h00006FA0 : data <= 8'b00000000 ;
			15'h00006FA1 : data <= 8'b00000000 ;
			15'h00006FA2 : data <= 8'b00000000 ;
			15'h00006FA3 : data <= 8'b00000000 ;
			15'h00006FA4 : data <= 8'b00000000 ;
			15'h00006FA5 : data <= 8'b00000000 ;
			15'h00006FA6 : data <= 8'b00000000 ;
			15'h00006FA7 : data <= 8'b00000000 ;
			15'h00006FA8 : data <= 8'b00000000 ;
			15'h00006FA9 : data <= 8'b00000000 ;
			15'h00006FAA : data <= 8'b00000000 ;
			15'h00006FAB : data <= 8'b00000000 ;
			15'h00006FAC : data <= 8'b00000000 ;
			15'h00006FAD : data <= 8'b00000000 ;
			15'h00006FAE : data <= 8'b00000000 ;
			15'h00006FAF : data <= 8'b00000000 ;
			15'h00006FB0 : data <= 8'b00000000 ;
			15'h00006FB1 : data <= 8'b00000000 ;
			15'h00006FB2 : data <= 8'b00000000 ;
			15'h00006FB3 : data <= 8'b00000000 ;
			15'h00006FB4 : data <= 8'b00000000 ;
			15'h00006FB5 : data <= 8'b00000000 ;
			15'h00006FB6 : data <= 8'b00000000 ;
			15'h00006FB7 : data <= 8'b00000000 ;
			15'h00006FB8 : data <= 8'b00000000 ;
			15'h00006FB9 : data <= 8'b00000000 ;
			15'h00006FBA : data <= 8'b00000000 ;
			15'h00006FBB : data <= 8'b00000000 ;
			15'h00006FBC : data <= 8'b00000000 ;
			15'h00006FBD : data <= 8'b00000000 ;
			15'h00006FBE : data <= 8'b00000000 ;
			15'h00006FBF : data <= 8'b00000000 ;
			15'h00006FC0 : data <= 8'b00000000 ;
			15'h00006FC1 : data <= 8'b00000000 ;
			15'h00006FC2 : data <= 8'b00000000 ;
			15'h00006FC3 : data <= 8'b00000000 ;
			15'h00006FC4 : data <= 8'b00000000 ;
			15'h00006FC5 : data <= 8'b00000000 ;
			15'h00006FC6 : data <= 8'b00000000 ;
			15'h00006FC7 : data <= 8'b00000000 ;
			15'h00006FC8 : data <= 8'b00000000 ;
			15'h00006FC9 : data <= 8'b00000000 ;
			15'h00006FCA : data <= 8'b00000000 ;
			15'h00006FCB : data <= 8'b00000000 ;
			15'h00006FCC : data <= 8'b00000000 ;
			15'h00006FCD : data <= 8'b00000000 ;
			15'h00006FCE : data <= 8'b00000000 ;
			15'h00006FCF : data <= 8'b00000000 ;
			15'h00006FD0 : data <= 8'b00000000 ;
			15'h00006FD1 : data <= 8'b00000000 ;
			15'h00006FD2 : data <= 8'b00000000 ;
			15'h00006FD3 : data <= 8'b00000000 ;
			15'h00006FD4 : data <= 8'b00000000 ;
			15'h00006FD5 : data <= 8'b00000000 ;
			15'h00006FD6 : data <= 8'b00000000 ;
			15'h00006FD7 : data <= 8'b00000000 ;
			15'h00006FD8 : data <= 8'b00000000 ;
			15'h00006FD9 : data <= 8'b00000000 ;
			15'h00006FDA : data <= 8'b00000000 ;
			15'h00006FDB : data <= 8'b00000000 ;
			15'h00006FDC : data <= 8'b00000000 ;
			15'h00006FDD : data <= 8'b00000000 ;
			15'h00006FDE : data <= 8'b00000000 ;
			15'h00006FDF : data <= 8'b00000000 ;
			15'h00006FE0 : data <= 8'b00000000 ;
			15'h00006FE1 : data <= 8'b00000000 ;
			15'h00006FE2 : data <= 8'b00000000 ;
			15'h00006FE3 : data <= 8'b00000000 ;
			15'h00006FE4 : data <= 8'b00000000 ;
			15'h00006FE5 : data <= 8'b00000000 ;
			15'h00006FE6 : data <= 8'b00000000 ;
			15'h00006FE7 : data <= 8'b00000000 ;
			15'h00006FE8 : data <= 8'b00000000 ;
			15'h00006FE9 : data <= 8'b00000000 ;
			15'h00006FEA : data <= 8'b00000000 ;
			15'h00006FEB : data <= 8'b00000000 ;
			15'h00006FEC : data <= 8'b00000000 ;
			15'h00006FED : data <= 8'b00000000 ;
			15'h00006FEE : data <= 8'b00000000 ;
			15'h00006FEF : data <= 8'b00000000 ;
			15'h00006FF0 : data <= 8'b00000000 ;
			15'h00006FF1 : data <= 8'b00000000 ;
			15'h00006FF2 : data <= 8'b00000000 ;
			15'h00006FF3 : data <= 8'b00000000 ;
			15'h00006FF4 : data <= 8'b00000000 ;
			15'h00006FF5 : data <= 8'b00000000 ;
			15'h00006FF6 : data <= 8'b00000000 ;
			15'h00006FF7 : data <= 8'b00000000 ;
			15'h00006FF8 : data <= 8'b00000000 ;
			15'h00006FF9 : data <= 8'b00000000 ;
			15'h00006FFA : data <= 8'b00000000 ;
			15'h00006FFB : data <= 8'b00000000 ;
			15'h00006FFC : data <= 8'b00000000 ;
			15'h00006FFD : data <= 8'b00000000 ;
			15'h00006FFE : data <= 8'b00000000 ;
			15'h00006FFF : data <= 8'b00000000 ;
			15'h00007000 : data <= 8'b00000000 ;
			15'h00007001 : data <= 8'b00000000 ;
			15'h00007002 : data <= 8'b00000000 ;
			15'h00007003 : data <= 8'b00000000 ;
			15'h00007004 : data <= 8'b00000000 ;
			15'h00007005 : data <= 8'b00000000 ;
			15'h00007006 : data <= 8'b00000000 ;
			15'h00007007 : data <= 8'b00000000 ;
			15'h00007008 : data <= 8'b00000000 ;
			15'h00007009 : data <= 8'b00000000 ;
			15'h0000700A : data <= 8'b00000000 ;
			15'h0000700B : data <= 8'b00000000 ;
			15'h0000700C : data <= 8'b00000000 ;
			15'h0000700D : data <= 8'b00000000 ;
			15'h0000700E : data <= 8'b00000000 ;
			15'h0000700F : data <= 8'b00000000 ;
			15'h00007010 : data <= 8'b00000000 ;
			15'h00007011 : data <= 8'b00000000 ;
			15'h00007012 : data <= 8'b00000000 ;
			15'h00007013 : data <= 8'b00000000 ;
			15'h00007014 : data <= 8'b00000000 ;
			15'h00007015 : data <= 8'b00000000 ;
			15'h00007016 : data <= 8'b00000000 ;
			15'h00007017 : data <= 8'b00000000 ;
			15'h00007018 : data <= 8'b00000000 ;
			15'h00007019 : data <= 8'b00000000 ;
			15'h0000701A : data <= 8'b00000000 ;
			15'h0000701B : data <= 8'b00000000 ;
			15'h0000701C : data <= 8'b00000000 ;
			15'h0000701D : data <= 8'b00000000 ;
			15'h0000701E : data <= 8'b00000000 ;
			15'h0000701F : data <= 8'b00000000 ;
			15'h00007020 : data <= 8'b00000000 ;
			15'h00007021 : data <= 8'b00000000 ;
			15'h00007022 : data <= 8'b00000000 ;
			15'h00007023 : data <= 8'b00000000 ;
			15'h00007024 : data <= 8'b00000000 ;
			15'h00007025 : data <= 8'b00000000 ;
			15'h00007026 : data <= 8'b00000000 ;
			15'h00007027 : data <= 8'b00000000 ;
			15'h00007028 : data <= 8'b00000000 ;
			15'h00007029 : data <= 8'b00000000 ;
			15'h0000702A : data <= 8'b00000000 ;
			15'h0000702B : data <= 8'b00000000 ;
			15'h0000702C : data <= 8'b00000000 ;
			15'h0000702D : data <= 8'b00000000 ;
			15'h0000702E : data <= 8'b00000000 ;
			15'h0000702F : data <= 8'b00000000 ;
			15'h00007030 : data <= 8'b00000000 ;
			15'h00007031 : data <= 8'b00000000 ;
			15'h00007032 : data <= 8'b00000000 ;
			15'h00007033 : data <= 8'b00000000 ;
			15'h00007034 : data <= 8'b00000000 ;
			15'h00007035 : data <= 8'b00000000 ;
			15'h00007036 : data <= 8'b00000000 ;
			15'h00007037 : data <= 8'b00000000 ;
			15'h00007038 : data <= 8'b00000000 ;
			15'h00007039 : data <= 8'b00000000 ;
			15'h0000703A : data <= 8'b00000000 ;
			15'h0000703B : data <= 8'b00000000 ;
			15'h0000703C : data <= 8'b00000000 ;
			15'h0000703D : data <= 8'b00000000 ;
			15'h0000703E : data <= 8'b00000000 ;
			15'h0000703F : data <= 8'b00000000 ;
			15'h00007040 : data <= 8'b00000000 ;
			15'h00007041 : data <= 8'b00000000 ;
			15'h00007042 : data <= 8'b00000000 ;
			15'h00007043 : data <= 8'b00000000 ;
			15'h00007044 : data <= 8'b00000000 ;
			15'h00007045 : data <= 8'b00000000 ;
			15'h00007046 : data <= 8'b00000000 ;
			15'h00007047 : data <= 8'b00000000 ;
			15'h00007048 : data <= 8'b00000000 ;
			15'h00007049 : data <= 8'b00000000 ;
			15'h0000704A : data <= 8'b00000000 ;
			15'h0000704B : data <= 8'b00000000 ;
			15'h0000704C : data <= 8'b00000000 ;
			15'h0000704D : data <= 8'b00000000 ;
			15'h0000704E : data <= 8'b00000000 ;
			15'h0000704F : data <= 8'b00000000 ;
			15'h00007050 : data <= 8'b00000000 ;
			15'h00007051 : data <= 8'b00000000 ;
			15'h00007052 : data <= 8'b00000000 ;
			15'h00007053 : data <= 8'b00000000 ;
			15'h00007054 : data <= 8'b00000000 ;
			15'h00007055 : data <= 8'b00000000 ;
			15'h00007056 : data <= 8'b00000000 ;
			15'h00007057 : data <= 8'b00000000 ;
			15'h00007058 : data <= 8'b00000000 ;
			15'h00007059 : data <= 8'b00000000 ;
			15'h0000705A : data <= 8'b00000000 ;
			15'h0000705B : data <= 8'b00000000 ;
			15'h0000705C : data <= 8'b00000000 ;
			15'h0000705D : data <= 8'b00000000 ;
			15'h0000705E : data <= 8'b00000000 ;
			15'h0000705F : data <= 8'b00000000 ;
			15'h00007060 : data <= 8'b00000000 ;
			15'h00007061 : data <= 8'b00000000 ;
			15'h00007062 : data <= 8'b00000000 ;
			15'h00007063 : data <= 8'b00000000 ;
			15'h00007064 : data <= 8'b00000000 ;
			15'h00007065 : data <= 8'b00000000 ;
			15'h00007066 : data <= 8'b00000000 ;
			15'h00007067 : data <= 8'b00000000 ;
			15'h00007068 : data <= 8'b00000000 ;
			15'h00007069 : data <= 8'b00000000 ;
			15'h0000706A : data <= 8'b00000000 ;
			15'h0000706B : data <= 8'b00000000 ;
			15'h0000706C : data <= 8'b00000000 ;
			15'h0000706D : data <= 8'b00000000 ;
			15'h0000706E : data <= 8'b00000000 ;
			15'h0000706F : data <= 8'b00000000 ;
			15'h00007070 : data <= 8'b00000000 ;
			15'h00007071 : data <= 8'b00000000 ;
			15'h00007072 : data <= 8'b00000000 ;
			15'h00007073 : data <= 8'b00000000 ;
			15'h00007074 : data <= 8'b00000000 ;
			15'h00007075 : data <= 8'b00000000 ;
			15'h00007076 : data <= 8'b00000000 ;
			15'h00007077 : data <= 8'b00000000 ;
			15'h00007078 : data <= 8'b00000000 ;
			15'h00007079 : data <= 8'b00000000 ;
			15'h0000707A : data <= 8'b00000000 ;
			15'h0000707B : data <= 8'b00000000 ;
			15'h0000707C : data <= 8'b00000000 ;
			15'h0000707D : data <= 8'b00000000 ;
			15'h0000707E : data <= 8'b00000000 ;
			15'h0000707F : data <= 8'b00000000 ;
			15'h00007080 : data <= 8'b00000000 ;
			15'h00007081 : data <= 8'b00000000 ;
			15'h00007082 : data <= 8'b00000000 ;
			15'h00007083 : data <= 8'b00000000 ;
			15'h00007084 : data <= 8'b00000000 ;
			15'h00007085 : data <= 8'b00000000 ;
			15'h00007086 : data <= 8'b00000000 ;
			15'h00007087 : data <= 8'b00000000 ;
			15'h00007088 : data <= 8'b00000000 ;
			15'h00007089 : data <= 8'b00000000 ;
			15'h0000708A : data <= 8'b00000000 ;
			15'h0000708B : data <= 8'b00000000 ;
			15'h0000708C : data <= 8'b00000000 ;
			15'h0000708D : data <= 8'b00000000 ;
			15'h0000708E : data <= 8'b00000000 ;
			15'h0000708F : data <= 8'b00000000 ;
			15'h00007090 : data <= 8'b00000000 ;
			15'h00007091 : data <= 8'b00000000 ;
			15'h00007092 : data <= 8'b00000000 ;
			15'h00007093 : data <= 8'b00000000 ;
			15'h00007094 : data <= 8'b00000000 ;
			15'h00007095 : data <= 8'b00000000 ;
			15'h00007096 : data <= 8'b00000000 ;
			15'h00007097 : data <= 8'b00000000 ;
			15'h00007098 : data <= 8'b00000000 ;
			15'h00007099 : data <= 8'b00000000 ;
			15'h0000709A : data <= 8'b00000000 ;
			15'h0000709B : data <= 8'b00000000 ;
			15'h0000709C : data <= 8'b00000000 ;
			15'h0000709D : data <= 8'b00000000 ;
			15'h0000709E : data <= 8'b00000000 ;
			15'h0000709F : data <= 8'b00000000 ;
			15'h000070A0 : data <= 8'b00000000 ;
			15'h000070A1 : data <= 8'b00000000 ;
			15'h000070A2 : data <= 8'b00000000 ;
			15'h000070A3 : data <= 8'b00000000 ;
			15'h000070A4 : data <= 8'b00000000 ;
			15'h000070A5 : data <= 8'b00000000 ;
			15'h000070A6 : data <= 8'b00000000 ;
			15'h000070A7 : data <= 8'b00000000 ;
			15'h000070A8 : data <= 8'b00000000 ;
			15'h000070A9 : data <= 8'b00000000 ;
			15'h000070AA : data <= 8'b00000000 ;
			15'h000070AB : data <= 8'b00000000 ;
			15'h000070AC : data <= 8'b00000000 ;
			15'h000070AD : data <= 8'b00000000 ;
			15'h000070AE : data <= 8'b00000000 ;
			15'h000070AF : data <= 8'b00000000 ;
			15'h000070B0 : data <= 8'b00000000 ;
			15'h000070B1 : data <= 8'b00000000 ;
			15'h000070B2 : data <= 8'b00000000 ;
			15'h000070B3 : data <= 8'b00000000 ;
			15'h000070B4 : data <= 8'b00000000 ;
			15'h000070B5 : data <= 8'b00000000 ;
			15'h000070B6 : data <= 8'b00000000 ;
			15'h000070B7 : data <= 8'b00000000 ;
			15'h000070B8 : data <= 8'b00000000 ;
			15'h000070B9 : data <= 8'b00000000 ;
			15'h000070BA : data <= 8'b00000000 ;
			15'h000070BB : data <= 8'b00000000 ;
			15'h000070BC : data <= 8'b00000000 ;
			15'h000070BD : data <= 8'b00000000 ;
			15'h000070BE : data <= 8'b00000000 ;
			15'h000070BF : data <= 8'b00000000 ;
			15'h000070C0 : data <= 8'b00000000 ;
			15'h000070C1 : data <= 8'b00000000 ;
			15'h000070C2 : data <= 8'b00000000 ;
			15'h000070C3 : data <= 8'b00000000 ;
			15'h000070C4 : data <= 8'b00000000 ;
			15'h000070C5 : data <= 8'b00000000 ;
			15'h000070C6 : data <= 8'b00000000 ;
			15'h000070C7 : data <= 8'b00000000 ;
			15'h000070C8 : data <= 8'b00000000 ;
			15'h000070C9 : data <= 8'b00000000 ;
			15'h000070CA : data <= 8'b00000000 ;
			15'h000070CB : data <= 8'b00000000 ;
			15'h000070CC : data <= 8'b00000000 ;
			15'h000070CD : data <= 8'b00000000 ;
			15'h000070CE : data <= 8'b00000000 ;
			15'h000070CF : data <= 8'b00000000 ;
			15'h000070D0 : data <= 8'b00000000 ;
			15'h000070D1 : data <= 8'b00000000 ;
			15'h000070D2 : data <= 8'b00000000 ;
			15'h000070D3 : data <= 8'b00000000 ;
			15'h000070D4 : data <= 8'b00000000 ;
			15'h000070D5 : data <= 8'b00000000 ;
			15'h000070D6 : data <= 8'b00000000 ;
			15'h000070D7 : data <= 8'b00000000 ;
			15'h000070D8 : data <= 8'b00000000 ;
			15'h000070D9 : data <= 8'b00000000 ;
			15'h000070DA : data <= 8'b00000000 ;
			15'h000070DB : data <= 8'b00000000 ;
			15'h000070DC : data <= 8'b00000000 ;
			15'h000070DD : data <= 8'b00000000 ;
			15'h000070DE : data <= 8'b00000000 ;
			15'h000070DF : data <= 8'b00000000 ;
			15'h000070E0 : data <= 8'b00000000 ;
			15'h000070E1 : data <= 8'b00000000 ;
			15'h000070E2 : data <= 8'b00000000 ;
			15'h000070E3 : data <= 8'b00000000 ;
			15'h000070E4 : data <= 8'b00000000 ;
			15'h000070E5 : data <= 8'b00000000 ;
			15'h000070E6 : data <= 8'b00000000 ;
			15'h000070E7 : data <= 8'b00000000 ;
			15'h000070E8 : data <= 8'b00000000 ;
			15'h000070E9 : data <= 8'b00000000 ;
			15'h000070EA : data <= 8'b00000000 ;
			15'h000070EB : data <= 8'b00000000 ;
			15'h000070EC : data <= 8'b00000000 ;
			15'h000070ED : data <= 8'b00000000 ;
			15'h000070EE : data <= 8'b00000000 ;
			15'h000070EF : data <= 8'b00000000 ;
			15'h000070F0 : data <= 8'b00000000 ;
			15'h000070F1 : data <= 8'b00000000 ;
			15'h000070F2 : data <= 8'b00000000 ;
			15'h000070F3 : data <= 8'b00000000 ;
			15'h000070F4 : data <= 8'b00000000 ;
			15'h000070F5 : data <= 8'b00000000 ;
			15'h000070F6 : data <= 8'b00000000 ;
			15'h000070F7 : data <= 8'b00000000 ;
			15'h000070F8 : data <= 8'b00000000 ;
			15'h000070F9 : data <= 8'b00000000 ;
			15'h000070FA : data <= 8'b00000000 ;
			15'h000070FB : data <= 8'b00000000 ;
			15'h000070FC : data <= 8'b00000000 ;
			15'h000070FD : data <= 8'b00000000 ;
			15'h000070FE : data <= 8'b00000000 ;
			15'h000070FF : data <= 8'b00000000 ;
			15'h00007100 : data <= 8'b00000000 ;
			15'h00007101 : data <= 8'b00000000 ;
			15'h00007102 : data <= 8'b00000000 ;
			15'h00007103 : data <= 8'b00000000 ;
			15'h00007104 : data <= 8'b00000000 ;
			15'h00007105 : data <= 8'b00000000 ;
			15'h00007106 : data <= 8'b00000000 ;
			15'h00007107 : data <= 8'b00000000 ;
			15'h00007108 : data <= 8'b00000000 ;
			15'h00007109 : data <= 8'b00000000 ;
			15'h0000710A : data <= 8'b00000000 ;
			15'h0000710B : data <= 8'b00000000 ;
			15'h0000710C : data <= 8'b00000000 ;
			15'h0000710D : data <= 8'b00000000 ;
			15'h0000710E : data <= 8'b00000000 ;
			15'h0000710F : data <= 8'b00000000 ;
			15'h00007110 : data <= 8'b00000000 ;
			15'h00007111 : data <= 8'b00000000 ;
			15'h00007112 : data <= 8'b00000000 ;
			15'h00007113 : data <= 8'b00000000 ;
			15'h00007114 : data <= 8'b00000000 ;
			15'h00007115 : data <= 8'b00000000 ;
			15'h00007116 : data <= 8'b00000000 ;
			15'h00007117 : data <= 8'b00000000 ;
			15'h00007118 : data <= 8'b00000000 ;
			15'h00007119 : data <= 8'b00000000 ;
			15'h0000711A : data <= 8'b00000000 ;
			15'h0000711B : data <= 8'b00000000 ;
			15'h0000711C : data <= 8'b00000000 ;
			15'h0000711D : data <= 8'b00000000 ;
			15'h0000711E : data <= 8'b00000000 ;
			15'h0000711F : data <= 8'b00000000 ;
			15'h00007120 : data <= 8'b00000000 ;
			15'h00007121 : data <= 8'b00000000 ;
			15'h00007122 : data <= 8'b00000000 ;
			15'h00007123 : data <= 8'b00000000 ;
			15'h00007124 : data <= 8'b00000000 ;
			15'h00007125 : data <= 8'b00000000 ;
			15'h00007126 : data <= 8'b00000000 ;
			15'h00007127 : data <= 8'b00000000 ;
			15'h00007128 : data <= 8'b00000000 ;
			15'h00007129 : data <= 8'b00000000 ;
			15'h0000712A : data <= 8'b00000000 ;
			15'h0000712B : data <= 8'b00000000 ;
			15'h0000712C : data <= 8'b00000000 ;
			15'h0000712D : data <= 8'b00000000 ;
			15'h0000712E : data <= 8'b00000000 ;
			15'h0000712F : data <= 8'b00000000 ;
			15'h00007130 : data <= 8'b00000000 ;
			15'h00007131 : data <= 8'b00000000 ;
			15'h00007132 : data <= 8'b00000000 ;
			15'h00007133 : data <= 8'b00000000 ;
			15'h00007134 : data <= 8'b00000000 ;
			15'h00007135 : data <= 8'b00000000 ;
			15'h00007136 : data <= 8'b00000000 ;
			15'h00007137 : data <= 8'b00000000 ;
			15'h00007138 : data <= 8'b00000000 ;
			15'h00007139 : data <= 8'b00000000 ;
			15'h0000713A : data <= 8'b00000000 ;
			15'h0000713B : data <= 8'b00000000 ;
			15'h0000713C : data <= 8'b00000000 ;
			15'h0000713D : data <= 8'b00000000 ;
			15'h0000713E : data <= 8'b00000000 ;
			15'h0000713F : data <= 8'b00000000 ;
			15'h00007140 : data <= 8'b00000000 ;
			15'h00007141 : data <= 8'b00000000 ;
			15'h00007142 : data <= 8'b00000000 ;
			15'h00007143 : data <= 8'b00000000 ;
			15'h00007144 : data <= 8'b00000000 ;
			15'h00007145 : data <= 8'b00000000 ;
			15'h00007146 : data <= 8'b00000000 ;
			15'h00007147 : data <= 8'b00000000 ;
			15'h00007148 : data <= 8'b00000000 ;
			15'h00007149 : data <= 8'b00000000 ;
			15'h0000714A : data <= 8'b00000000 ;
			15'h0000714B : data <= 8'b00000000 ;
			15'h0000714C : data <= 8'b00000000 ;
			15'h0000714D : data <= 8'b00000000 ;
			15'h0000714E : data <= 8'b00000000 ;
			15'h0000714F : data <= 8'b00000000 ;
			15'h00007150 : data <= 8'b00000000 ;
			15'h00007151 : data <= 8'b00000000 ;
			15'h00007152 : data <= 8'b00000000 ;
			15'h00007153 : data <= 8'b00000000 ;
			15'h00007154 : data <= 8'b00000000 ;
			15'h00007155 : data <= 8'b00000000 ;
			15'h00007156 : data <= 8'b00000000 ;
			15'h00007157 : data <= 8'b00000000 ;
			15'h00007158 : data <= 8'b00000000 ;
			15'h00007159 : data <= 8'b00000000 ;
			15'h0000715A : data <= 8'b00000000 ;
			15'h0000715B : data <= 8'b00000000 ;
			15'h0000715C : data <= 8'b00000000 ;
			15'h0000715D : data <= 8'b00000000 ;
			15'h0000715E : data <= 8'b00000000 ;
			15'h0000715F : data <= 8'b00000000 ;
			15'h00007160 : data <= 8'b00000000 ;
			15'h00007161 : data <= 8'b00000000 ;
			15'h00007162 : data <= 8'b00000000 ;
			15'h00007163 : data <= 8'b00000000 ;
			15'h00007164 : data <= 8'b00000000 ;
			15'h00007165 : data <= 8'b00000000 ;
			15'h00007166 : data <= 8'b00000000 ;
			15'h00007167 : data <= 8'b00000000 ;
			15'h00007168 : data <= 8'b00000000 ;
			15'h00007169 : data <= 8'b00000000 ;
			15'h0000716A : data <= 8'b00000000 ;
			15'h0000716B : data <= 8'b00000000 ;
			15'h0000716C : data <= 8'b00000000 ;
			15'h0000716D : data <= 8'b00000000 ;
			15'h0000716E : data <= 8'b00000000 ;
			15'h0000716F : data <= 8'b00000000 ;
			15'h00007170 : data <= 8'b00000000 ;
			15'h00007171 : data <= 8'b00000000 ;
			15'h00007172 : data <= 8'b00000000 ;
			15'h00007173 : data <= 8'b00000000 ;
			15'h00007174 : data <= 8'b00000000 ;
			15'h00007175 : data <= 8'b00000000 ;
			15'h00007176 : data <= 8'b00000000 ;
			15'h00007177 : data <= 8'b00000000 ;
			15'h00007178 : data <= 8'b00000000 ;
			15'h00007179 : data <= 8'b00000000 ;
			15'h0000717A : data <= 8'b00000000 ;
			15'h0000717B : data <= 8'b00000000 ;
			15'h0000717C : data <= 8'b00000000 ;
			15'h0000717D : data <= 8'b00000000 ;
			15'h0000717E : data <= 8'b00000000 ;
			15'h0000717F : data <= 8'b00000000 ;
			15'h00007180 : data <= 8'b00000000 ;
			15'h00007181 : data <= 8'b00000000 ;
			15'h00007182 : data <= 8'b00000000 ;
			15'h00007183 : data <= 8'b00000000 ;
			15'h00007184 : data <= 8'b00000000 ;
			15'h00007185 : data <= 8'b00000000 ;
			15'h00007186 : data <= 8'b00000000 ;
			15'h00007187 : data <= 8'b00000000 ;
			15'h00007188 : data <= 8'b00000000 ;
			15'h00007189 : data <= 8'b00000000 ;
			15'h0000718A : data <= 8'b00000000 ;
			15'h0000718B : data <= 8'b00000000 ;
			15'h0000718C : data <= 8'b00000000 ;
			15'h0000718D : data <= 8'b00000000 ;
			15'h0000718E : data <= 8'b00000000 ;
			15'h0000718F : data <= 8'b00000000 ;
			15'h00007190 : data <= 8'b00000000 ;
			15'h00007191 : data <= 8'b00000000 ;
			15'h00007192 : data <= 8'b00000000 ;
			15'h00007193 : data <= 8'b00000000 ;
			15'h00007194 : data <= 8'b00000000 ;
			15'h00007195 : data <= 8'b00000000 ;
			15'h00007196 : data <= 8'b00000000 ;
			15'h00007197 : data <= 8'b00000000 ;
			15'h00007198 : data <= 8'b00000000 ;
			15'h00007199 : data <= 8'b00000000 ;
			15'h0000719A : data <= 8'b00000000 ;
			15'h0000719B : data <= 8'b00000000 ;
			15'h0000719C : data <= 8'b00000000 ;
			15'h0000719D : data <= 8'b00000000 ;
			15'h0000719E : data <= 8'b00000000 ;
			15'h0000719F : data <= 8'b00000000 ;
			15'h000071A0 : data <= 8'b00000000 ;
			15'h000071A1 : data <= 8'b00000000 ;
			15'h000071A2 : data <= 8'b00000000 ;
			15'h000071A3 : data <= 8'b00000000 ;
			15'h000071A4 : data <= 8'b00000000 ;
			15'h000071A5 : data <= 8'b00000000 ;
			15'h000071A6 : data <= 8'b00000000 ;
			15'h000071A7 : data <= 8'b00000000 ;
			15'h000071A8 : data <= 8'b00000000 ;
			15'h000071A9 : data <= 8'b00000000 ;
			15'h000071AA : data <= 8'b00000000 ;
			15'h000071AB : data <= 8'b00000000 ;
			15'h000071AC : data <= 8'b00000000 ;
			15'h000071AD : data <= 8'b00000000 ;
			15'h000071AE : data <= 8'b00000000 ;
			15'h000071AF : data <= 8'b00000000 ;
			15'h000071B0 : data <= 8'b00000000 ;
			15'h000071B1 : data <= 8'b00000000 ;
			15'h000071B2 : data <= 8'b00000000 ;
			15'h000071B3 : data <= 8'b00000000 ;
			15'h000071B4 : data <= 8'b00000000 ;
			15'h000071B5 : data <= 8'b00000000 ;
			15'h000071B6 : data <= 8'b00000000 ;
			15'h000071B7 : data <= 8'b00000000 ;
			15'h000071B8 : data <= 8'b00000000 ;
			15'h000071B9 : data <= 8'b00000000 ;
			15'h000071BA : data <= 8'b00000000 ;
			15'h000071BB : data <= 8'b00000000 ;
			15'h000071BC : data <= 8'b00000000 ;
			15'h000071BD : data <= 8'b00000000 ;
			15'h000071BE : data <= 8'b00000000 ;
			15'h000071BF : data <= 8'b00000000 ;
			15'h000071C0 : data <= 8'b00000000 ;
			15'h000071C1 : data <= 8'b00000000 ;
			15'h000071C2 : data <= 8'b00000000 ;
			15'h000071C3 : data <= 8'b00000000 ;
			15'h000071C4 : data <= 8'b00000000 ;
			15'h000071C5 : data <= 8'b00000000 ;
			15'h000071C6 : data <= 8'b00000000 ;
			15'h000071C7 : data <= 8'b00000000 ;
			15'h000071C8 : data <= 8'b00000000 ;
			15'h000071C9 : data <= 8'b00000000 ;
			15'h000071CA : data <= 8'b00000000 ;
			15'h000071CB : data <= 8'b00000000 ;
			15'h000071CC : data <= 8'b00000000 ;
			15'h000071CD : data <= 8'b00000000 ;
			15'h000071CE : data <= 8'b00000000 ;
			15'h000071CF : data <= 8'b00000000 ;
			15'h000071D0 : data <= 8'b00000000 ;
			15'h000071D1 : data <= 8'b00000000 ;
			15'h000071D2 : data <= 8'b00000000 ;
			15'h000071D3 : data <= 8'b00000000 ;
			15'h000071D4 : data <= 8'b00000000 ;
			15'h000071D5 : data <= 8'b00000000 ;
			15'h000071D6 : data <= 8'b00000000 ;
			15'h000071D7 : data <= 8'b00000000 ;
			15'h000071D8 : data <= 8'b00000000 ;
			15'h000071D9 : data <= 8'b00000000 ;
			15'h000071DA : data <= 8'b00000000 ;
			15'h000071DB : data <= 8'b00000000 ;
			15'h000071DC : data <= 8'b00000000 ;
			15'h000071DD : data <= 8'b00000000 ;
			15'h000071DE : data <= 8'b00000000 ;
			15'h000071DF : data <= 8'b00000000 ;
			15'h000071E0 : data <= 8'b00000000 ;
			15'h000071E1 : data <= 8'b00000000 ;
			15'h000071E2 : data <= 8'b00000000 ;
			15'h000071E3 : data <= 8'b00000000 ;
			15'h000071E4 : data <= 8'b00000000 ;
			15'h000071E5 : data <= 8'b00000000 ;
			15'h000071E6 : data <= 8'b00000000 ;
			15'h000071E7 : data <= 8'b00000000 ;
			15'h000071E8 : data <= 8'b00000000 ;
			15'h000071E9 : data <= 8'b00000000 ;
			15'h000071EA : data <= 8'b00000000 ;
			15'h000071EB : data <= 8'b00000000 ;
			15'h000071EC : data <= 8'b00000000 ;
			15'h000071ED : data <= 8'b00000000 ;
			15'h000071EE : data <= 8'b00000000 ;
			15'h000071EF : data <= 8'b00000000 ;
			15'h000071F0 : data <= 8'b00000000 ;
			15'h000071F1 : data <= 8'b00000000 ;
			15'h000071F2 : data <= 8'b00000000 ;
			15'h000071F3 : data <= 8'b00000000 ;
			15'h000071F4 : data <= 8'b00000000 ;
			15'h000071F5 : data <= 8'b00000000 ;
			15'h000071F6 : data <= 8'b00000000 ;
			15'h000071F7 : data <= 8'b00000000 ;
			15'h000071F8 : data <= 8'b00000000 ;
			15'h000071F9 : data <= 8'b00000000 ;
			15'h000071FA : data <= 8'b00000000 ;
			15'h000071FB : data <= 8'b00000000 ;
			15'h000071FC : data <= 8'b00000000 ;
			15'h000071FD : data <= 8'b00000000 ;
			15'h000071FE : data <= 8'b00000000 ;
			15'h000071FF : data <= 8'b00000000 ;
			15'h00007200 : data <= 8'b00000000 ;
			15'h00007201 : data <= 8'b00000000 ;
			15'h00007202 : data <= 8'b00000000 ;
			15'h00007203 : data <= 8'b00000000 ;
			15'h00007204 : data <= 8'b00000000 ;
			15'h00007205 : data <= 8'b00000000 ;
			15'h00007206 : data <= 8'b00000000 ;
			15'h00007207 : data <= 8'b00000000 ;
			15'h00007208 : data <= 8'b00000000 ;
			15'h00007209 : data <= 8'b00000000 ;
			15'h0000720A : data <= 8'b00000000 ;
			15'h0000720B : data <= 8'b00000000 ;
			15'h0000720C : data <= 8'b00000000 ;
			15'h0000720D : data <= 8'b00000000 ;
			15'h0000720E : data <= 8'b00000000 ;
			15'h0000720F : data <= 8'b00000000 ;
			15'h00007210 : data <= 8'b00000000 ;
			15'h00007211 : data <= 8'b00000000 ;
			15'h00007212 : data <= 8'b00000000 ;
			15'h00007213 : data <= 8'b00000000 ;
			15'h00007214 : data <= 8'b00000000 ;
			15'h00007215 : data <= 8'b00000000 ;
			15'h00007216 : data <= 8'b00000000 ;
			15'h00007217 : data <= 8'b00000000 ;
			15'h00007218 : data <= 8'b00000000 ;
			15'h00007219 : data <= 8'b00000000 ;
			15'h0000721A : data <= 8'b00000000 ;
			15'h0000721B : data <= 8'b00000000 ;
			15'h0000721C : data <= 8'b00000000 ;
			15'h0000721D : data <= 8'b00000000 ;
			15'h0000721E : data <= 8'b00000000 ;
			15'h0000721F : data <= 8'b00000000 ;
			15'h00007220 : data <= 8'b00000000 ;
			15'h00007221 : data <= 8'b00000000 ;
			15'h00007222 : data <= 8'b00000000 ;
			15'h00007223 : data <= 8'b00000000 ;
			15'h00007224 : data <= 8'b00000000 ;
			15'h00007225 : data <= 8'b00000000 ;
			15'h00007226 : data <= 8'b00000000 ;
			15'h00007227 : data <= 8'b00000000 ;
			15'h00007228 : data <= 8'b00000000 ;
			15'h00007229 : data <= 8'b00000000 ;
			15'h0000722A : data <= 8'b00000000 ;
			15'h0000722B : data <= 8'b00000000 ;
			15'h0000722C : data <= 8'b00000000 ;
			15'h0000722D : data <= 8'b00000000 ;
			15'h0000722E : data <= 8'b00000000 ;
			15'h0000722F : data <= 8'b00000000 ;
			15'h00007230 : data <= 8'b00000000 ;
			15'h00007231 : data <= 8'b00000000 ;
			15'h00007232 : data <= 8'b00000000 ;
			15'h00007233 : data <= 8'b00000000 ;
			15'h00007234 : data <= 8'b00000000 ;
			15'h00007235 : data <= 8'b00000000 ;
			15'h00007236 : data <= 8'b00000000 ;
			15'h00007237 : data <= 8'b00000000 ;
			15'h00007238 : data <= 8'b00000000 ;
			15'h00007239 : data <= 8'b00000000 ;
			15'h0000723A : data <= 8'b00000000 ;
			15'h0000723B : data <= 8'b00000000 ;
			15'h0000723C : data <= 8'b00000000 ;
			15'h0000723D : data <= 8'b00000000 ;
			15'h0000723E : data <= 8'b00000000 ;
			15'h0000723F : data <= 8'b00000000 ;
			15'h00007240 : data <= 8'b00000000 ;
			15'h00007241 : data <= 8'b00000000 ;
			15'h00007242 : data <= 8'b00000000 ;
			15'h00007243 : data <= 8'b00000000 ;
			15'h00007244 : data <= 8'b00000000 ;
			15'h00007245 : data <= 8'b00000000 ;
			15'h00007246 : data <= 8'b00000000 ;
			15'h00007247 : data <= 8'b00000000 ;
			15'h00007248 : data <= 8'b00000000 ;
			15'h00007249 : data <= 8'b00000000 ;
			15'h0000724A : data <= 8'b00000000 ;
			15'h0000724B : data <= 8'b00000000 ;
			15'h0000724C : data <= 8'b00000000 ;
			15'h0000724D : data <= 8'b00000000 ;
			15'h0000724E : data <= 8'b00000000 ;
			15'h0000724F : data <= 8'b00000000 ;
			15'h00007250 : data <= 8'b00000000 ;
			15'h00007251 : data <= 8'b00000000 ;
			15'h00007252 : data <= 8'b00000000 ;
			15'h00007253 : data <= 8'b00000000 ;
			15'h00007254 : data <= 8'b00000000 ;
			15'h00007255 : data <= 8'b00000000 ;
			15'h00007256 : data <= 8'b00000000 ;
			15'h00007257 : data <= 8'b00000000 ;
			15'h00007258 : data <= 8'b00000000 ;
			15'h00007259 : data <= 8'b00000000 ;
			15'h0000725A : data <= 8'b00000000 ;
			15'h0000725B : data <= 8'b00000000 ;
			15'h0000725C : data <= 8'b00000000 ;
			15'h0000725D : data <= 8'b00000000 ;
			15'h0000725E : data <= 8'b00000000 ;
			15'h0000725F : data <= 8'b00000000 ;
			15'h00007260 : data <= 8'b00000000 ;
			15'h00007261 : data <= 8'b00000000 ;
			15'h00007262 : data <= 8'b00000000 ;
			15'h00007263 : data <= 8'b00000000 ;
			15'h00007264 : data <= 8'b00000000 ;
			15'h00007265 : data <= 8'b00000000 ;
			15'h00007266 : data <= 8'b00000000 ;
			15'h00007267 : data <= 8'b00000000 ;
			15'h00007268 : data <= 8'b00000000 ;
			15'h00007269 : data <= 8'b00000000 ;
			15'h0000726A : data <= 8'b00000000 ;
			15'h0000726B : data <= 8'b00000000 ;
			15'h0000726C : data <= 8'b00000000 ;
			15'h0000726D : data <= 8'b00000000 ;
			15'h0000726E : data <= 8'b00000000 ;
			15'h0000726F : data <= 8'b00000000 ;
			15'h00007270 : data <= 8'b00000000 ;
			15'h00007271 : data <= 8'b00000000 ;
			15'h00007272 : data <= 8'b00000000 ;
			15'h00007273 : data <= 8'b00000000 ;
			15'h00007274 : data <= 8'b00000000 ;
			15'h00007275 : data <= 8'b00000000 ;
			15'h00007276 : data <= 8'b00000000 ;
			15'h00007277 : data <= 8'b00000000 ;
			15'h00007278 : data <= 8'b00000000 ;
			15'h00007279 : data <= 8'b00000000 ;
			15'h0000727A : data <= 8'b00000000 ;
			15'h0000727B : data <= 8'b00000000 ;
			15'h0000727C : data <= 8'b00000000 ;
			15'h0000727D : data <= 8'b00000000 ;
			15'h0000727E : data <= 8'b00000000 ;
			15'h0000727F : data <= 8'b00000000 ;
			15'h00007280 : data <= 8'b00000000 ;
			15'h00007281 : data <= 8'b00000000 ;
			15'h00007282 : data <= 8'b00000000 ;
			15'h00007283 : data <= 8'b00000000 ;
			15'h00007284 : data <= 8'b00000000 ;
			15'h00007285 : data <= 8'b00000000 ;
			15'h00007286 : data <= 8'b00000000 ;
			15'h00007287 : data <= 8'b00000000 ;
			15'h00007288 : data <= 8'b00000000 ;
			15'h00007289 : data <= 8'b00000000 ;
			15'h0000728A : data <= 8'b00000000 ;
			15'h0000728B : data <= 8'b00000000 ;
			15'h0000728C : data <= 8'b00000000 ;
			15'h0000728D : data <= 8'b00000000 ;
			15'h0000728E : data <= 8'b00000000 ;
			15'h0000728F : data <= 8'b00000000 ;
			15'h00007290 : data <= 8'b00000000 ;
			15'h00007291 : data <= 8'b00000000 ;
			15'h00007292 : data <= 8'b00000000 ;
			15'h00007293 : data <= 8'b00000000 ;
			15'h00007294 : data <= 8'b00000000 ;
			15'h00007295 : data <= 8'b00000000 ;
			15'h00007296 : data <= 8'b00000000 ;
			15'h00007297 : data <= 8'b00000000 ;
			15'h00007298 : data <= 8'b00000000 ;
			15'h00007299 : data <= 8'b00000000 ;
			15'h0000729A : data <= 8'b00000000 ;
			15'h0000729B : data <= 8'b00000000 ;
			15'h0000729C : data <= 8'b00000000 ;
			15'h0000729D : data <= 8'b00000000 ;
			15'h0000729E : data <= 8'b00000000 ;
			15'h0000729F : data <= 8'b00000000 ;
			15'h000072A0 : data <= 8'b00000000 ;
			15'h000072A1 : data <= 8'b00000000 ;
			15'h000072A2 : data <= 8'b00000000 ;
			15'h000072A3 : data <= 8'b00000000 ;
			15'h000072A4 : data <= 8'b00000000 ;
			15'h000072A5 : data <= 8'b00000000 ;
			15'h000072A6 : data <= 8'b00000000 ;
			15'h000072A7 : data <= 8'b00000000 ;
			15'h000072A8 : data <= 8'b00000000 ;
			15'h000072A9 : data <= 8'b00000000 ;
			15'h000072AA : data <= 8'b00000000 ;
			15'h000072AB : data <= 8'b00000000 ;
			15'h000072AC : data <= 8'b00000000 ;
			15'h000072AD : data <= 8'b00000000 ;
			15'h000072AE : data <= 8'b00000000 ;
			15'h000072AF : data <= 8'b00000000 ;
			15'h000072B0 : data <= 8'b00000000 ;
			15'h000072B1 : data <= 8'b00000000 ;
			15'h000072B2 : data <= 8'b00000000 ;
			15'h000072B3 : data <= 8'b00000000 ;
			15'h000072B4 : data <= 8'b00000000 ;
			15'h000072B5 : data <= 8'b00000000 ;
			15'h000072B6 : data <= 8'b00000000 ;
			15'h000072B7 : data <= 8'b00000000 ;
			15'h000072B8 : data <= 8'b00000000 ;
			15'h000072B9 : data <= 8'b00000000 ;
			15'h000072BA : data <= 8'b00000000 ;
			15'h000072BB : data <= 8'b00000000 ;
			15'h000072BC : data <= 8'b00000000 ;
			15'h000072BD : data <= 8'b00000000 ;
			15'h000072BE : data <= 8'b00000000 ;
			15'h000072BF : data <= 8'b00000000 ;
			15'h000072C0 : data <= 8'b00000000 ;
			15'h000072C1 : data <= 8'b00000000 ;
			15'h000072C2 : data <= 8'b00000000 ;
			15'h000072C3 : data <= 8'b00000000 ;
			15'h000072C4 : data <= 8'b00000000 ;
			15'h000072C5 : data <= 8'b00000000 ;
			15'h000072C6 : data <= 8'b00000000 ;
			15'h000072C7 : data <= 8'b00000000 ;
			15'h000072C8 : data <= 8'b00000000 ;
			15'h000072C9 : data <= 8'b00000000 ;
			15'h000072CA : data <= 8'b00000000 ;
			15'h000072CB : data <= 8'b00000000 ;
			15'h000072CC : data <= 8'b00000000 ;
			15'h000072CD : data <= 8'b00000000 ;
			15'h000072CE : data <= 8'b00000000 ;
			15'h000072CF : data <= 8'b00000000 ;
			15'h000072D0 : data <= 8'b00000000 ;
			15'h000072D1 : data <= 8'b00000000 ;
			15'h000072D2 : data <= 8'b00000000 ;
			15'h000072D3 : data <= 8'b00000000 ;
			15'h000072D4 : data <= 8'b00000000 ;
			15'h000072D5 : data <= 8'b00000000 ;
			15'h000072D6 : data <= 8'b00000000 ;
			15'h000072D7 : data <= 8'b00000000 ;
			15'h000072D8 : data <= 8'b00000000 ;
			15'h000072D9 : data <= 8'b00000000 ;
			15'h000072DA : data <= 8'b00000000 ;
			15'h000072DB : data <= 8'b00000000 ;
			15'h000072DC : data <= 8'b00000000 ;
			15'h000072DD : data <= 8'b00000000 ;
			15'h000072DE : data <= 8'b00000000 ;
			15'h000072DF : data <= 8'b00000000 ;
			15'h000072E0 : data <= 8'b00000000 ;
			15'h000072E1 : data <= 8'b00000000 ;
			15'h000072E2 : data <= 8'b00000000 ;
			15'h000072E3 : data <= 8'b00000000 ;
			15'h000072E4 : data <= 8'b00000000 ;
			15'h000072E5 : data <= 8'b00000000 ;
			15'h000072E6 : data <= 8'b00000000 ;
			15'h000072E7 : data <= 8'b00000000 ;
			15'h000072E8 : data <= 8'b00000000 ;
			15'h000072E9 : data <= 8'b00000000 ;
			15'h000072EA : data <= 8'b00000000 ;
			15'h000072EB : data <= 8'b00000000 ;
			15'h000072EC : data <= 8'b00000000 ;
			15'h000072ED : data <= 8'b00000000 ;
			15'h000072EE : data <= 8'b00000000 ;
			15'h000072EF : data <= 8'b00000000 ;
			15'h000072F0 : data <= 8'b00000000 ;
			15'h000072F1 : data <= 8'b00000000 ;
			15'h000072F2 : data <= 8'b00000000 ;
			15'h000072F3 : data <= 8'b00000000 ;
			15'h000072F4 : data <= 8'b00000000 ;
			15'h000072F5 : data <= 8'b00000000 ;
			15'h000072F6 : data <= 8'b00000000 ;
			15'h000072F7 : data <= 8'b00000000 ;
			15'h000072F8 : data <= 8'b00000000 ;
			15'h000072F9 : data <= 8'b00000000 ;
			15'h000072FA : data <= 8'b00000000 ;
			15'h000072FB : data <= 8'b00000000 ;
			15'h000072FC : data <= 8'b00000000 ;
			15'h000072FD : data <= 8'b00000000 ;
			15'h000072FE : data <= 8'b00000000 ;
			15'h000072FF : data <= 8'b00000000 ;
			15'h00007300 : data <= 8'b00000000 ;
			15'h00007301 : data <= 8'b00000000 ;
			15'h00007302 : data <= 8'b00000000 ;
			15'h00007303 : data <= 8'b00000000 ;
			15'h00007304 : data <= 8'b00000000 ;
			15'h00007305 : data <= 8'b00000000 ;
			15'h00007306 : data <= 8'b00000000 ;
			15'h00007307 : data <= 8'b00000000 ;
			15'h00007308 : data <= 8'b00000000 ;
			15'h00007309 : data <= 8'b00000000 ;
			15'h0000730A : data <= 8'b00000000 ;
			15'h0000730B : data <= 8'b00000000 ;
			15'h0000730C : data <= 8'b00000000 ;
			15'h0000730D : data <= 8'b00000000 ;
			15'h0000730E : data <= 8'b00000000 ;
			15'h0000730F : data <= 8'b00000000 ;
			15'h00007310 : data <= 8'b00000000 ;
			15'h00007311 : data <= 8'b00000000 ;
			15'h00007312 : data <= 8'b00000000 ;
			15'h00007313 : data <= 8'b00000000 ;
			15'h00007314 : data <= 8'b00000000 ;
			15'h00007315 : data <= 8'b00000000 ;
			15'h00007316 : data <= 8'b00000000 ;
			15'h00007317 : data <= 8'b00000000 ;
			15'h00007318 : data <= 8'b00000000 ;
			15'h00007319 : data <= 8'b00000000 ;
			15'h0000731A : data <= 8'b00000000 ;
			15'h0000731B : data <= 8'b00000000 ;
			15'h0000731C : data <= 8'b00000000 ;
			15'h0000731D : data <= 8'b00000000 ;
			15'h0000731E : data <= 8'b00000000 ;
			15'h0000731F : data <= 8'b00000000 ;
			15'h00007320 : data <= 8'b00000000 ;
			15'h00007321 : data <= 8'b00000000 ;
			15'h00007322 : data <= 8'b00000000 ;
			15'h00007323 : data <= 8'b00000000 ;
			15'h00007324 : data <= 8'b00000000 ;
			15'h00007325 : data <= 8'b00000000 ;
			15'h00007326 : data <= 8'b00000000 ;
			15'h00007327 : data <= 8'b00000000 ;
			15'h00007328 : data <= 8'b00000000 ;
			15'h00007329 : data <= 8'b00000000 ;
			15'h0000732A : data <= 8'b00000000 ;
			15'h0000732B : data <= 8'b00000000 ;
			15'h0000732C : data <= 8'b00000000 ;
			15'h0000732D : data <= 8'b00000000 ;
			15'h0000732E : data <= 8'b00000000 ;
			15'h0000732F : data <= 8'b00000000 ;
			15'h00007330 : data <= 8'b00000000 ;
			15'h00007331 : data <= 8'b00000000 ;
			15'h00007332 : data <= 8'b00000000 ;
			15'h00007333 : data <= 8'b00000000 ;
			15'h00007334 : data <= 8'b00000000 ;
			15'h00007335 : data <= 8'b00000000 ;
			15'h00007336 : data <= 8'b00000000 ;
			15'h00007337 : data <= 8'b00000000 ;
			15'h00007338 : data <= 8'b00000000 ;
			15'h00007339 : data <= 8'b00000000 ;
			15'h0000733A : data <= 8'b00000000 ;
			15'h0000733B : data <= 8'b00000000 ;
			15'h0000733C : data <= 8'b00000000 ;
			15'h0000733D : data <= 8'b00000000 ;
			15'h0000733E : data <= 8'b00000000 ;
			15'h0000733F : data <= 8'b00000000 ;
			15'h00007340 : data <= 8'b00000000 ;
			15'h00007341 : data <= 8'b00000000 ;
			15'h00007342 : data <= 8'b00000000 ;
			15'h00007343 : data <= 8'b00000000 ;
			15'h00007344 : data <= 8'b00000000 ;
			15'h00007345 : data <= 8'b00000000 ;
			15'h00007346 : data <= 8'b00000000 ;
			15'h00007347 : data <= 8'b00000000 ;
			15'h00007348 : data <= 8'b00000000 ;
			15'h00007349 : data <= 8'b00000000 ;
			15'h0000734A : data <= 8'b00000000 ;
			15'h0000734B : data <= 8'b00000000 ;
			15'h0000734C : data <= 8'b00000000 ;
			15'h0000734D : data <= 8'b00000000 ;
			15'h0000734E : data <= 8'b00000000 ;
			15'h0000734F : data <= 8'b00000000 ;
			15'h00007350 : data <= 8'b00000000 ;
			15'h00007351 : data <= 8'b00000000 ;
			15'h00007352 : data <= 8'b00000000 ;
			15'h00007353 : data <= 8'b00000000 ;
			15'h00007354 : data <= 8'b00000000 ;
			15'h00007355 : data <= 8'b00000000 ;
			15'h00007356 : data <= 8'b00000000 ;
			15'h00007357 : data <= 8'b00000000 ;
			15'h00007358 : data <= 8'b00000000 ;
			15'h00007359 : data <= 8'b00000000 ;
			15'h0000735A : data <= 8'b00000000 ;
			15'h0000735B : data <= 8'b00000000 ;
			15'h0000735C : data <= 8'b00000000 ;
			15'h0000735D : data <= 8'b00000000 ;
			15'h0000735E : data <= 8'b00000000 ;
			15'h0000735F : data <= 8'b00000000 ;
			15'h00007360 : data <= 8'b00000000 ;
			15'h00007361 : data <= 8'b00000000 ;
			15'h00007362 : data <= 8'b00000000 ;
			15'h00007363 : data <= 8'b00000000 ;
			15'h00007364 : data <= 8'b00000000 ;
			15'h00007365 : data <= 8'b00000000 ;
			15'h00007366 : data <= 8'b00000000 ;
			15'h00007367 : data <= 8'b00000000 ;
			15'h00007368 : data <= 8'b00000000 ;
			15'h00007369 : data <= 8'b00000000 ;
			15'h0000736A : data <= 8'b00000000 ;
			15'h0000736B : data <= 8'b00000000 ;
			15'h0000736C : data <= 8'b00000000 ;
			15'h0000736D : data <= 8'b00000000 ;
			15'h0000736E : data <= 8'b00000000 ;
			15'h0000736F : data <= 8'b00000000 ;
			15'h00007370 : data <= 8'b00000000 ;
			15'h00007371 : data <= 8'b00000000 ;
			15'h00007372 : data <= 8'b00000000 ;
			15'h00007373 : data <= 8'b00000000 ;
			15'h00007374 : data <= 8'b00000000 ;
			15'h00007375 : data <= 8'b00000000 ;
			15'h00007376 : data <= 8'b00000000 ;
			15'h00007377 : data <= 8'b00000000 ;
			15'h00007378 : data <= 8'b00000000 ;
			15'h00007379 : data <= 8'b00000000 ;
			15'h0000737A : data <= 8'b00000000 ;
			15'h0000737B : data <= 8'b00000000 ;
			15'h0000737C : data <= 8'b00000000 ;
			15'h0000737D : data <= 8'b00000000 ;
			15'h0000737E : data <= 8'b00000000 ;
			15'h0000737F : data <= 8'b00000000 ;
			15'h00007380 : data <= 8'b00000000 ;
			15'h00007381 : data <= 8'b00000000 ;
			15'h00007382 : data <= 8'b00000000 ;
			15'h00007383 : data <= 8'b00000000 ;
			15'h00007384 : data <= 8'b00000000 ;
			15'h00007385 : data <= 8'b00000000 ;
			15'h00007386 : data <= 8'b00000000 ;
			15'h00007387 : data <= 8'b00000000 ;
			15'h00007388 : data <= 8'b00000000 ;
			15'h00007389 : data <= 8'b00000000 ;
			15'h0000738A : data <= 8'b00000000 ;
			15'h0000738B : data <= 8'b00000000 ;
			15'h0000738C : data <= 8'b00000000 ;
			15'h0000738D : data <= 8'b00000000 ;
			15'h0000738E : data <= 8'b00000000 ;
			15'h0000738F : data <= 8'b00000000 ;
			15'h00007390 : data <= 8'b00000000 ;
			15'h00007391 : data <= 8'b00000000 ;
			15'h00007392 : data <= 8'b00000000 ;
			15'h00007393 : data <= 8'b00000000 ;
			15'h00007394 : data <= 8'b00000000 ;
			15'h00007395 : data <= 8'b00000000 ;
			15'h00007396 : data <= 8'b00000000 ;
			15'h00007397 : data <= 8'b00000000 ;
			15'h00007398 : data <= 8'b00000000 ;
			15'h00007399 : data <= 8'b00000000 ;
			15'h0000739A : data <= 8'b00000000 ;
			15'h0000739B : data <= 8'b00000000 ;
			15'h0000739C : data <= 8'b00000000 ;
			15'h0000739D : data <= 8'b00000000 ;
			15'h0000739E : data <= 8'b00000000 ;
			15'h0000739F : data <= 8'b00000000 ;
			15'h000073A0 : data <= 8'b00000000 ;
			15'h000073A1 : data <= 8'b00000000 ;
			15'h000073A2 : data <= 8'b00000000 ;
			15'h000073A3 : data <= 8'b00000000 ;
			15'h000073A4 : data <= 8'b00000000 ;
			15'h000073A5 : data <= 8'b00000000 ;
			15'h000073A6 : data <= 8'b00000000 ;
			15'h000073A7 : data <= 8'b00000000 ;
			15'h000073A8 : data <= 8'b00000000 ;
			15'h000073A9 : data <= 8'b00000000 ;
			15'h000073AA : data <= 8'b00000000 ;
			15'h000073AB : data <= 8'b00000000 ;
			15'h000073AC : data <= 8'b00000000 ;
			15'h000073AD : data <= 8'b00000000 ;
			15'h000073AE : data <= 8'b00000000 ;
			15'h000073AF : data <= 8'b00000000 ;
			15'h000073B0 : data <= 8'b00000000 ;
			15'h000073B1 : data <= 8'b00000000 ;
			15'h000073B2 : data <= 8'b00000000 ;
			15'h000073B3 : data <= 8'b00000000 ;
			15'h000073B4 : data <= 8'b00000000 ;
			15'h000073B5 : data <= 8'b00000000 ;
			15'h000073B6 : data <= 8'b00000000 ;
			15'h000073B7 : data <= 8'b00000000 ;
			15'h000073B8 : data <= 8'b00000000 ;
			15'h000073B9 : data <= 8'b00000000 ;
			15'h000073BA : data <= 8'b00000000 ;
			15'h000073BB : data <= 8'b00000000 ;
			15'h000073BC : data <= 8'b00000000 ;
			15'h000073BD : data <= 8'b00000000 ;
			15'h000073BE : data <= 8'b00000000 ;
			15'h000073BF : data <= 8'b00000000 ;
			15'h000073C0 : data <= 8'b00000000 ;
			15'h000073C1 : data <= 8'b00000000 ;
			15'h000073C2 : data <= 8'b00000000 ;
			15'h000073C3 : data <= 8'b00000000 ;
			15'h000073C4 : data <= 8'b00000000 ;
			15'h000073C5 : data <= 8'b00000000 ;
			15'h000073C6 : data <= 8'b00000000 ;
			15'h000073C7 : data <= 8'b00000000 ;
			15'h000073C8 : data <= 8'b00000000 ;
			15'h000073C9 : data <= 8'b00000000 ;
			15'h000073CA : data <= 8'b00000000 ;
			15'h000073CB : data <= 8'b00000000 ;
			15'h000073CC : data <= 8'b00000000 ;
			15'h000073CD : data <= 8'b00000000 ;
			15'h000073CE : data <= 8'b00000000 ;
			15'h000073CF : data <= 8'b00000000 ;
			15'h000073D0 : data <= 8'b00000000 ;
			15'h000073D1 : data <= 8'b00000000 ;
			15'h000073D2 : data <= 8'b00000000 ;
			15'h000073D3 : data <= 8'b00000000 ;
			15'h000073D4 : data <= 8'b00000000 ;
			15'h000073D5 : data <= 8'b00000000 ;
			15'h000073D6 : data <= 8'b00000000 ;
			15'h000073D7 : data <= 8'b00000000 ;
			15'h000073D8 : data <= 8'b00000000 ;
			15'h000073D9 : data <= 8'b00000000 ;
			15'h000073DA : data <= 8'b00000000 ;
			15'h000073DB : data <= 8'b00000000 ;
			15'h000073DC : data <= 8'b00000000 ;
			15'h000073DD : data <= 8'b00000000 ;
			15'h000073DE : data <= 8'b00000000 ;
			15'h000073DF : data <= 8'b00000000 ;
			15'h000073E0 : data <= 8'b00000000 ;
			15'h000073E1 : data <= 8'b00000000 ;
			15'h000073E2 : data <= 8'b00000000 ;
			15'h000073E3 : data <= 8'b00000000 ;
			15'h000073E4 : data <= 8'b00000000 ;
			15'h000073E5 : data <= 8'b00000000 ;
			15'h000073E6 : data <= 8'b00000000 ;
			15'h000073E7 : data <= 8'b00000000 ;
			15'h000073E8 : data <= 8'b00000000 ;
			15'h000073E9 : data <= 8'b00000000 ;
			15'h000073EA : data <= 8'b00000000 ;
			15'h000073EB : data <= 8'b00000000 ;
			15'h000073EC : data <= 8'b00000000 ;
			15'h000073ED : data <= 8'b00000000 ;
			15'h000073EE : data <= 8'b00000000 ;
			15'h000073EF : data <= 8'b00000000 ;
			15'h000073F0 : data <= 8'b00000000 ;
			15'h000073F1 : data <= 8'b00000000 ;
			15'h000073F2 : data <= 8'b00000000 ;
			15'h000073F3 : data <= 8'b00000000 ;
			15'h000073F4 : data <= 8'b00000000 ;
			15'h000073F5 : data <= 8'b00000000 ;
			15'h000073F6 : data <= 8'b00000000 ;
			15'h000073F7 : data <= 8'b00000000 ;
			15'h000073F8 : data <= 8'b00000000 ;
			15'h000073F9 : data <= 8'b00000000 ;
			15'h000073FA : data <= 8'b00000000 ;
			15'h000073FB : data <= 8'b00000000 ;
			15'h000073FC : data <= 8'b00000000 ;
			15'h000073FD : data <= 8'b00000000 ;
			15'h000073FE : data <= 8'b00000000 ;
			15'h000073FF : data <= 8'b00000000 ;
			15'h00007400 : data <= 8'b00000000 ;
			15'h00007401 : data <= 8'b00000000 ;
			15'h00007402 : data <= 8'b00000000 ;
			15'h00007403 : data <= 8'b00000000 ;
			15'h00007404 : data <= 8'b00000000 ;
			15'h00007405 : data <= 8'b00000000 ;
			15'h00007406 : data <= 8'b00000000 ;
			15'h00007407 : data <= 8'b00000000 ;
			15'h00007408 : data <= 8'b00000000 ;
			15'h00007409 : data <= 8'b00000000 ;
			15'h0000740A : data <= 8'b00000000 ;
			15'h0000740B : data <= 8'b00000000 ;
			15'h0000740C : data <= 8'b00000000 ;
			15'h0000740D : data <= 8'b00000000 ;
			15'h0000740E : data <= 8'b00000000 ;
			15'h0000740F : data <= 8'b00000000 ;
			15'h00007410 : data <= 8'b00000000 ;
			15'h00007411 : data <= 8'b00000000 ;
			15'h00007412 : data <= 8'b00000000 ;
			15'h00007413 : data <= 8'b00000000 ;
			15'h00007414 : data <= 8'b00000000 ;
			15'h00007415 : data <= 8'b00000000 ;
			15'h00007416 : data <= 8'b00000000 ;
			15'h00007417 : data <= 8'b00000000 ;
			15'h00007418 : data <= 8'b00000000 ;
			15'h00007419 : data <= 8'b00000000 ;
			15'h0000741A : data <= 8'b00000000 ;
			15'h0000741B : data <= 8'b00000000 ;
			15'h0000741C : data <= 8'b00000000 ;
			15'h0000741D : data <= 8'b00000000 ;
			15'h0000741E : data <= 8'b00000000 ;
			15'h0000741F : data <= 8'b00000000 ;
			15'h00007420 : data <= 8'b00000000 ;
			15'h00007421 : data <= 8'b00000000 ;
			15'h00007422 : data <= 8'b00000000 ;
			15'h00007423 : data <= 8'b00000000 ;
			15'h00007424 : data <= 8'b00000000 ;
			15'h00007425 : data <= 8'b00000000 ;
			15'h00007426 : data <= 8'b00000000 ;
			15'h00007427 : data <= 8'b00000000 ;
			15'h00007428 : data <= 8'b00000000 ;
			15'h00007429 : data <= 8'b00000000 ;
			15'h0000742A : data <= 8'b00000000 ;
			15'h0000742B : data <= 8'b00000000 ;
			15'h0000742C : data <= 8'b00000000 ;
			15'h0000742D : data <= 8'b00000000 ;
			15'h0000742E : data <= 8'b00000000 ;
			15'h0000742F : data <= 8'b00000000 ;
			15'h00007430 : data <= 8'b00000000 ;
			15'h00007431 : data <= 8'b00000000 ;
			15'h00007432 : data <= 8'b00000000 ;
			15'h00007433 : data <= 8'b00000000 ;
			15'h00007434 : data <= 8'b00000000 ;
			15'h00007435 : data <= 8'b00000000 ;
			15'h00007436 : data <= 8'b00000000 ;
			15'h00007437 : data <= 8'b00000000 ;
			15'h00007438 : data <= 8'b00000000 ;
			15'h00007439 : data <= 8'b00000000 ;
			15'h0000743A : data <= 8'b00000000 ;
			15'h0000743B : data <= 8'b00000000 ;
			15'h0000743C : data <= 8'b00000000 ;
			15'h0000743D : data <= 8'b00000000 ;
			15'h0000743E : data <= 8'b00000000 ;
			15'h0000743F : data <= 8'b00000000 ;
			15'h00007440 : data <= 8'b00000000 ;
			15'h00007441 : data <= 8'b00000000 ;
			15'h00007442 : data <= 8'b00000000 ;
			15'h00007443 : data <= 8'b00000000 ;
			15'h00007444 : data <= 8'b00000000 ;
			15'h00007445 : data <= 8'b00000000 ;
			15'h00007446 : data <= 8'b00000000 ;
			15'h00007447 : data <= 8'b00000000 ;
			15'h00007448 : data <= 8'b00000000 ;
			15'h00007449 : data <= 8'b00000000 ;
			15'h0000744A : data <= 8'b00000000 ;
			15'h0000744B : data <= 8'b00000000 ;
			15'h0000744C : data <= 8'b00000000 ;
			15'h0000744D : data <= 8'b00000000 ;
			15'h0000744E : data <= 8'b00000000 ;
			15'h0000744F : data <= 8'b00000000 ;
			15'h00007450 : data <= 8'b00000000 ;
			15'h00007451 : data <= 8'b00000000 ;
			15'h00007452 : data <= 8'b00000000 ;
			15'h00007453 : data <= 8'b00000000 ;
			15'h00007454 : data <= 8'b00000000 ;
			15'h00007455 : data <= 8'b00000000 ;
			15'h00007456 : data <= 8'b00000000 ;
			15'h00007457 : data <= 8'b00000000 ;
			15'h00007458 : data <= 8'b00000000 ;
			15'h00007459 : data <= 8'b00000000 ;
			15'h0000745A : data <= 8'b00000000 ;
			15'h0000745B : data <= 8'b00000000 ;
			15'h0000745C : data <= 8'b00000000 ;
			15'h0000745D : data <= 8'b00000000 ;
			15'h0000745E : data <= 8'b00000000 ;
			15'h0000745F : data <= 8'b00000000 ;
			15'h00007460 : data <= 8'b00000000 ;
			15'h00007461 : data <= 8'b00000000 ;
			15'h00007462 : data <= 8'b00000000 ;
			15'h00007463 : data <= 8'b00000000 ;
			15'h00007464 : data <= 8'b00000000 ;
			15'h00007465 : data <= 8'b00000000 ;
			15'h00007466 : data <= 8'b00000000 ;
			15'h00007467 : data <= 8'b00000000 ;
			15'h00007468 : data <= 8'b00000000 ;
			15'h00007469 : data <= 8'b00000000 ;
			15'h0000746A : data <= 8'b00000000 ;
			15'h0000746B : data <= 8'b00000000 ;
			15'h0000746C : data <= 8'b00000000 ;
			15'h0000746D : data <= 8'b00000000 ;
			15'h0000746E : data <= 8'b00000000 ;
			15'h0000746F : data <= 8'b00000000 ;
			15'h00007470 : data <= 8'b00000000 ;
			15'h00007471 : data <= 8'b00000000 ;
			15'h00007472 : data <= 8'b00000000 ;
			15'h00007473 : data <= 8'b00000000 ;
			15'h00007474 : data <= 8'b00000000 ;
			15'h00007475 : data <= 8'b00000000 ;
			15'h00007476 : data <= 8'b00000000 ;
			15'h00007477 : data <= 8'b00000000 ;
			15'h00007478 : data <= 8'b00000000 ;
			15'h00007479 : data <= 8'b00000000 ;
			15'h0000747A : data <= 8'b00000000 ;
			15'h0000747B : data <= 8'b00000000 ;
			15'h0000747C : data <= 8'b00000000 ;
			15'h0000747D : data <= 8'b00000000 ;
			15'h0000747E : data <= 8'b00000000 ;
			15'h0000747F : data <= 8'b00000000 ;
			15'h00007480 : data <= 8'b00000000 ;
			15'h00007481 : data <= 8'b00000000 ;
			15'h00007482 : data <= 8'b00000000 ;
			15'h00007483 : data <= 8'b00000000 ;
			15'h00007484 : data <= 8'b00000000 ;
			15'h00007485 : data <= 8'b00000000 ;
			15'h00007486 : data <= 8'b00000000 ;
			15'h00007487 : data <= 8'b00000000 ;
			15'h00007488 : data <= 8'b00000000 ;
			15'h00007489 : data <= 8'b00000000 ;
			15'h0000748A : data <= 8'b00000000 ;
			15'h0000748B : data <= 8'b00000000 ;
			15'h0000748C : data <= 8'b00000000 ;
			15'h0000748D : data <= 8'b00000000 ;
			15'h0000748E : data <= 8'b00000000 ;
			15'h0000748F : data <= 8'b00000000 ;
			15'h00007490 : data <= 8'b00000000 ;
			15'h00007491 : data <= 8'b00000000 ;
			15'h00007492 : data <= 8'b00000000 ;
			15'h00007493 : data <= 8'b00000000 ;
			15'h00007494 : data <= 8'b00000000 ;
			15'h00007495 : data <= 8'b00000000 ;
			15'h00007496 : data <= 8'b00000000 ;
			15'h00007497 : data <= 8'b00000000 ;
			15'h00007498 : data <= 8'b00000000 ;
			15'h00007499 : data <= 8'b00000000 ;
			15'h0000749A : data <= 8'b00000000 ;
			15'h0000749B : data <= 8'b00000000 ;
			15'h0000749C : data <= 8'b00000000 ;
			15'h0000749D : data <= 8'b00000000 ;
			15'h0000749E : data <= 8'b00000000 ;
			15'h0000749F : data <= 8'b00000000 ;
			15'h000074A0 : data <= 8'b00000000 ;
			15'h000074A1 : data <= 8'b00000000 ;
			15'h000074A2 : data <= 8'b00000000 ;
			15'h000074A3 : data <= 8'b00000000 ;
			15'h000074A4 : data <= 8'b00000000 ;
			15'h000074A5 : data <= 8'b00000000 ;
			15'h000074A6 : data <= 8'b00000000 ;
			15'h000074A7 : data <= 8'b00000000 ;
			15'h000074A8 : data <= 8'b00000000 ;
			15'h000074A9 : data <= 8'b00000000 ;
			15'h000074AA : data <= 8'b00000000 ;
			15'h000074AB : data <= 8'b00000000 ;
			15'h000074AC : data <= 8'b00000000 ;
			15'h000074AD : data <= 8'b00000000 ;
			15'h000074AE : data <= 8'b00000000 ;
			15'h000074AF : data <= 8'b00000000 ;
			15'h000074B0 : data <= 8'b00000000 ;
			15'h000074B1 : data <= 8'b00000000 ;
			15'h000074B2 : data <= 8'b00000000 ;
			15'h000074B3 : data <= 8'b00000000 ;
			15'h000074B4 : data <= 8'b00000000 ;
			15'h000074B5 : data <= 8'b00000000 ;
			15'h000074B6 : data <= 8'b00000000 ;
			15'h000074B7 : data <= 8'b00000000 ;
			15'h000074B8 : data <= 8'b00000000 ;
			15'h000074B9 : data <= 8'b00000000 ;
			15'h000074BA : data <= 8'b00000000 ;
			15'h000074BB : data <= 8'b00000000 ;
			15'h000074BC : data <= 8'b00000000 ;
			15'h000074BD : data <= 8'b00000000 ;
			15'h000074BE : data <= 8'b00000000 ;
			15'h000074BF : data <= 8'b00000000 ;
			15'h000074C0 : data <= 8'b00000000 ;
			15'h000074C1 : data <= 8'b00000000 ;
			15'h000074C2 : data <= 8'b00000000 ;
			15'h000074C3 : data <= 8'b00000000 ;
			15'h000074C4 : data <= 8'b00000000 ;
			15'h000074C5 : data <= 8'b00000000 ;
			15'h000074C6 : data <= 8'b00000000 ;
			15'h000074C7 : data <= 8'b00000000 ;
			15'h000074C8 : data <= 8'b00000000 ;
			15'h000074C9 : data <= 8'b00000000 ;
			15'h000074CA : data <= 8'b00000000 ;
			15'h000074CB : data <= 8'b00000000 ;
			15'h000074CC : data <= 8'b00000000 ;
			15'h000074CD : data <= 8'b00000000 ;
			15'h000074CE : data <= 8'b00000000 ;
			15'h000074CF : data <= 8'b00000000 ;
			15'h000074D0 : data <= 8'b00000000 ;
			15'h000074D1 : data <= 8'b00000000 ;
			15'h000074D2 : data <= 8'b00000000 ;
			15'h000074D3 : data <= 8'b00000000 ;
			15'h000074D4 : data <= 8'b00000000 ;
			15'h000074D5 : data <= 8'b00000000 ;
			15'h000074D6 : data <= 8'b00000000 ;
			15'h000074D7 : data <= 8'b00000000 ;
			15'h000074D8 : data <= 8'b00000000 ;
			15'h000074D9 : data <= 8'b00000000 ;
			15'h000074DA : data <= 8'b00000000 ;
			15'h000074DB : data <= 8'b00000000 ;
			15'h000074DC : data <= 8'b00000000 ;
			15'h000074DD : data <= 8'b00000000 ;
			15'h000074DE : data <= 8'b00000000 ;
			15'h000074DF : data <= 8'b00000000 ;
			15'h000074E0 : data <= 8'b00000000 ;
			15'h000074E1 : data <= 8'b00000000 ;
			15'h000074E2 : data <= 8'b00000000 ;
			15'h000074E3 : data <= 8'b00000000 ;
			15'h000074E4 : data <= 8'b00000000 ;
			15'h000074E5 : data <= 8'b00000000 ;
			15'h000074E6 : data <= 8'b00000000 ;
			15'h000074E7 : data <= 8'b00000000 ;
			15'h000074E8 : data <= 8'b00000000 ;
			15'h000074E9 : data <= 8'b00000000 ;
			15'h000074EA : data <= 8'b00000000 ;
			15'h000074EB : data <= 8'b00000000 ;
			15'h000074EC : data <= 8'b00000000 ;
			15'h000074ED : data <= 8'b00000000 ;
			15'h000074EE : data <= 8'b00000000 ;
			15'h000074EF : data <= 8'b00000000 ;
			15'h000074F0 : data <= 8'b00000000 ;
			15'h000074F1 : data <= 8'b00000000 ;
			15'h000074F2 : data <= 8'b00000000 ;
			15'h000074F3 : data <= 8'b00000000 ;
			15'h000074F4 : data <= 8'b00000000 ;
			15'h000074F5 : data <= 8'b00000000 ;
			15'h000074F6 : data <= 8'b00000000 ;
			15'h000074F7 : data <= 8'b00000000 ;
			15'h000074F8 : data <= 8'b00000000 ;
			15'h000074F9 : data <= 8'b00000000 ;
			15'h000074FA : data <= 8'b00000000 ;
			15'h000074FB : data <= 8'b00000000 ;
			15'h000074FC : data <= 8'b00000000 ;
			15'h000074FD : data <= 8'b00000000 ;
			15'h000074FE : data <= 8'b00000000 ;
			15'h000074FF : data <= 8'b00000000 ;
			15'h00007500 : data <= 8'b00000000 ;
			15'h00007501 : data <= 8'b00000000 ;
			15'h00007502 : data <= 8'b00000000 ;
			15'h00007503 : data <= 8'b00000000 ;
			15'h00007504 : data <= 8'b00000000 ;
			15'h00007505 : data <= 8'b00000000 ;
			15'h00007506 : data <= 8'b00000000 ;
			15'h00007507 : data <= 8'b00000000 ;
			15'h00007508 : data <= 8'b00000000 ;
			15'h00007509 : data <= 8'b00000000 ;
			15'h0000750A : data <= 8'b00000000 ;
			15'h0000750B : data <= 8'b00000000 ;
			15'h0000750C : data <= 8'b00000000 ;
			15'h0000750D : data <= 8'b00000000 ;
			15'h0000750E : data <= 8'b00000000 ;
			15'h0000750F : data <= 8'b00000000 ;
			15'h00007510 : data <= 8'b00000000 ;
			15'h00007511 : data <= 8'b00000000 ;
			15'h00007512 : data <= 8'b00000000 ;
			15'h00007513 : data <= 8'b00000000 ;
			15'h00007514 : data <= 8'b00000000 ;
			15'h00007515 : data <= 8'b00000000 ;
			15'h00007516 : data <= 8'b00000000 ;
			15'h00007517 : data <= 8'b00000000 ;
			15'h00007518 : data <= 8'b00000000 ;
			15'h00007519 : data <= 8'b00000000 ;
			15'h0000751A : data <= 8'b00000000 ;
			15'h0000751B : data <= 8'b00000000 ;
			15'h0000751C : data <= 8'b00000000 ;
			15'h0000751D : data <= 8'b00000000 ;
			15'h0000751E : data <= 8'b00000000 ;
			15'h0000751F : data <= 8'b00000000 ;
			15'h00007520 : data <= 8'b00000000 ;
			15'h00007521 : data <= 8'b00000000 ;
			15'h00007522 : data <= 8'b00000000 ;
			15'h00007523 : data <= 8'b00000000 ;
			15'h00007524 : data <= 8'b00000000 ;
			15'h00007525 : data <= 8'b00000000 ;
			15'h00007526 : data <= 8'b00000000 ;
			15'h00007527 : data <= 8'b00000000 ;
			15'h00007528 : data <= 8'b00000000 ;
			15'h00007529 : data <= 8'b00000000 ;
			15'h0000752A : data <= 8'b00000000 ;
			15'h0000752B : data <= 8'b00000000 ;
			15'h0000752C : data <= 8'b00000000 ;
			15'h0000752D : data <= 8'b00000000 ;
			15'h0000752E : data <= 8'b00000000 ;
			15'h0000752F : data <= 8'b00000000 ;
			15'h00007530 : data <= 8'b00000000 ;
			15'h00007531 : data <= 8'b00000000 ;
			15'h00007532 : data <= 8'b00000000 ;
			15'h00007533 : data <= 8'b00000000 ;
			15'h00007534 : data <= 8'b00000000 ;
			15'h00007535 : data <= 8'b00000000 ;
			15'h00007536 : data <= 8'b00000000 ;
			15'h00007537 : data <= 8'b00000000 ;
			15'h00007538 : data <= 8'b00000000 ;
			15'h00007539 : data <= 8'b00000000 ;
			15'h0000753A : data <= 8'b00000000 ;
			15'h0000753B : data <= 8'b00000000 ;
			15'h0000753C : data <= 8'b00000000 ;
			15'h0000753D : data <= 8'b00000000 ;
			15'h0000753E : data <= 8'b00000000 ;
			15'h0000753F : data <= 8'b00000000 ;
			15'h00007540 : data <= 8'b00000000 ;
			15'h00007541 : data <= 8'b00000000 ;
			15'h00007542 : data <= 8'b00000000 ;
			15'h00007543 : data <= 8'b00000000 ;
			15'h00007544 : data <= 8'b00000000 ;
			15'h00007545 : data <= 8'b00000000 ;
			15'h00007546 : data <= 8'b00000000 ;
			15'h00007547 : data <= 8'b00000000 ;
			15'h00007548 : data <= 8'b00000000 ;
			15'h00007549 : data <= 8'b00000000 ;
			15'h0000754A : data <= 8'b00000000 ;
			15'h0000754B : data <= 8'b00000000 ;
			15'h0000754C : data <= 8'b00000000 ;
			15'h0000754D : data <= 8'b00000000 ;
			15'h0000754E : data <= 8'b00000000 ;
			15'h0000754F : data <= 8'b00000000 ;
			15'h00007550 : data <= 8'b00000000 ;
			15'h00007551 : data <= 8'b00000000 ;
			15'h00007552 : data <= 8'b00000000 ;
			15'h00007553 : data <= 8'b00000000 ;
			15'h00007554 : data <= 8'b00000000 ;
			15'h00007555 : data <= 8'b00000000 ;
			15'h00007556 : data <= 8'b00000000 ;
			15'h00007557 : data <= 8'b00000000 ;
			15'h00007558 : data <= 8'b00000000 ;
			15'h00007559 : data <= 8'b00000000 ;
			15'h0000755A : data <= 8'b00000000 ;
			15'h0000755B : data <= 8'b00000000 ;
			15'h0000755C : data <= 8'b00000000 ;
			15'h0000755D : data <= 8'b00000000 ;
			15'h0000755E : data <= 8'b00000000 ;
			15'h0000755F : data <= 8'b00000000 ;
			15'h00007560 : data <= 8'b00000000 ;
			15'h00007561 : data <= 8'b00000000 ;
			15'h00007562 : data <= 8'b00000000 ;
			15'h00007563 : data <= 8'b00000000 ;
			15'h00007564 : data <= 8'b00000000 ;
			15'h00007565 : data <= 8'b00000000 ;
			15'h00007566 : data <= 8'b00000000 ;
			15'h00007567 : data <= 8'b00000000 ;
			15'h00007568 : data <= 8'b00000000 ;
			15'h00007569 : data <= 8'b00000000 ;
			15'h0000756A : data <= 8'b00000000 ;
			15'h0000756B : data <= 8'b00000000 ;
			15'h0000756C : data <= 8'b00000000 ;
			15'h0000756D : data <= 8'b00000000 ;
			15'h0000756E : data <= 8'b00000000 ;
			15'h0000756F : data <= 8'b00000000 ;
			15'h00007570 : data <= 8'b00000000 ;
			15'h00007571 : data <= 8'b00000000 ;
			15'h00007572 : data <= 8'b00000000 ;
			15'h00007573 : data <= 8'b00000000 ;
			15'h00007574 : data <= 8'b00000000 ;
			15'h00007575 : data <= 8'b00000000 ;
			15'h00007576 : data <= 8'b00000000 ;
			15'h00007577 : data <= 8'b00000000 ;
			15'h00007578 : data <= 8'b00000000 ;
			15'h00007579 : data <= 8'b00000000 ;
			15'h0000757A : data <= 8'b00000000 ;
			15'h0000757B : data <= 8'b00000000 ;
			15'h0000757C : data <= 8'b00000000 ;
			15'h0000757D : data <= 8'b00000000 ;
			15'h0000757E : data <= 8'b00000000 ;
			15'h0000757F : data <= 8'b00000000 ;
			15'h00007580 : data <= 8'b00000000 ;
			15'h00007581 : data <= 8'b00000000 ;
			15'h00007582 : data <= 8'b00000000 ;
			15'h00007583 : data <= 8'b00000000 ;
			15'h00007584 : data <= 8'b00000000 ;
			15'h00007585 : data <= 8'b00000000 ;
			15'h00007586 : data <= 8'b00000000 ;
			15'h00007587 : data <= 8'b00000000 ;
			15'h00007588 : data <= 8'b00000000 ;
			15'h00007589 : data <= 8'b00000000 ;
			15'h0000758A : data <= 8'b00000000 ;
			15'h0000758B : data <= 8'b00000000 ;
			15'h0000758C : data <= 8'b00000000 ;
			15'h0000758D : data <= 8'b00000000 ;
			15'h0000758E : data <= 8'b00000000 ;
			15'h0000758F : data <= 8'b00000000 ;
			15'h00007590 : data <= 8'b00000000 ;
			15'h00007591 : data <= 8'b00000000 ;
			15'h00007592 : data <= 8'b00000000 ;
			15'h00007593 : data <= 8'b00000000 ;
			15'h00007594 : data <= 8'b00000000 ;
			15'h00007595 : data <= 8'b00000000 ;
			15'h00007596 : data <= 8'b00000000 ;
			15'h00007597 : data <= 8'b00000000 ;
			15'h00007598 : data <= 8'b00000000 ;
			15'h00007599 : data <= 8'b00000000 ;
			15'h0000759A : data <= 8'b00000000 ;
			15'h0000759B : data <= 8'b00000000 ;
			15'h0000759C : data <= 8'b00000000 ;
			15'h0000759D : data <= 8'b00000000 ;
			15'h0000759E : data <= 8'b00000000 ;
			15'h0000759F : data <= 8'b00000000 ;
			15'h000075A0 : data <= 8'b00000000 ;
			15'h000075A1 : data <= 8'b00000000 ;
			15'h000075A2 : data <= 8'b00000000 ;
			15'h000075A3 : data <= 8'b00000000 ;
			15'h000075A4 : data <= 8'b00000000 ;
			15'h000075A5 : data <= 8'b00000000 ;
			15'h000075A6 : data <= 8'b00000000 ;
			15'h000075A7 : data <= 8'b00000000 ;
			15'h000075A8 : data <= 8'b00000000 ;
			15'h000075A9 : data <= 8'b00000000 ;
			15'h000075AA : data <= 8'b00000000 ;
			15'h000075AB : data <= 8'b00000000 ;
			15'h000075AC : data <= 8'b00000000 ;
			15'h000075AD : data <= 8'b00000000 ;
			15'h000075AE : data <= 8'b00000000 ;
			15'h000075AF : data <= 8'b00000000 ;
			15'h000075B0 : data <= 8'b00000000 ;
			15'h000075B1 : data <= 8'b00000000 ;
			15'h000075B2 : data <= 8'b00000000 ;
			15'h000075B3 : data <= 8'b00000000 ;
			15'h000075B4 : data <= 8'b00000000 ;
			15'h000075B5 : data <= 8'b00000000 ;
			15'h000075B6 : data <= 8'b00000000 ;
			15'h000075B7 : data <= 8'b00000000 ;
			15'h000075B8 : data <= 8'b00000000 ;
			15'h000075B9 : data <= 8'b00000000 ;
			15'h000075BA : data <= 8'b00000000 ;
			15'h000075BB : data <= 8'b00000000 ;
			15'h000075BC : data <= 8'b00000000 ;
			15'h000075BD : data <= 8'b00000000 ;
			15'h000075BE : data <= 8'b00000000 ;
			15'h000075BF : data <= 8'b00000000 ;
			15'h000075C0 : data <= 8'b00000000 ;
			15'h000075C1 : data <= 8'b00000000 ;
			15'h000075C2 : data <= 8'b00000000 ;
			15'h000075C3 : data <= 8'b00000000 ;
			15'h000075C4 : data <= 8'b00000000 ;
			15'h000075C5 : data <= 8'b00000000 ;
			15'h000075C6 : data <= 8'b00000000 ;
			15'h000075C7 : data <= 8'b00000000 ;
			15'h000075C8 : data <= 8'b00000000 ;
			15'h000075C9 : data <= 8'b00000000 ;
			15'h000075CA : data <= 8'b00000000 ;
			15'h000075CB : data <= 8'b00000000 ;
			15'h000075CC : data <= 8'b00000000 ;
			15'h000075CD : data <= 8'b00000000 ;
			15'h000075CE : data <= 8'b00000000 ;
			15'h000075CF : data <= 8'b00000000 ;
			15'h000075D0 : data <= 8'b00000000 ;
			15'h000075D1 : data <= 8'b00000000 ;
			15'h000075D2 : data <= 8'b00000000 ;
			15'h000075D3 : data <= 8'b00000000 ;
			15'h000075D4 : data <= 8'b00000000 ;
			15'h000075D5 : data <= 8'b00000000 ;
			15'h000075D6 : data <= 8'b00000000 ;
			15'h000075D7 : data <= 8'b00000000 ;
			15'h000075D8 : data <= 8'b00000000 ;
			15'h000075D9 : data <= 8'b00000000 ;
			15'h000075DA : data <= 8'b00000000 ;
			15'h000075DB : data <= 8'b00000000 ;
			15'h000075DC : data <= 8'b00000000 ;
			15'h000075DD : data <= 8'b00000000 ;
			15'h000075DE : data <= 8'b00000000 ;
			15'h000075DF : data <= 8'b00000000 ;
			15'h000075E0 : data <= 8'b00000000 ;
			15'h000075E1 : data <= 8'b00000000 ;
			15'h000075E2 : data <= 8'b00000000 ;
			15'h000075E3 : data <= 8'b00000000 ;
			15'h000075E4 : data <= 8'b00000000 ;
			15'h000075E5 : data <= 8'b00000000 ;
			15'h000075E6 : data <= 8'b00000000 ;
			15'h000075E7 : data <= 8'b00000000 ;
			15'h000075E8 : data <= 8'b00000000 ;
			15'h000075E9 : data <= 8'b00000000 ;
			15'h000075EA : data <= 8'b00000000 ;
			15'h000075EB : data <= 8'b00000000 ;
			15'h000075EC : data <= 8'b00000000 ;
			15'h000075ED : data <= 8'b00000000 ;
			15'h000075EE : data <= 8'b00000000 ;
			15'h000075EF : data <= 8'b00000000 ;
			15'h000075F0 : data <= 8'b00000000 ;
			15'h000075F1 : data <= 8'b00000000 ;
			15'h000075F2 : data <= 8'b00000000 ;
			15'h000075F3 : data <= 8'b00000000 ;
			15'h000075F4 : data <= 8'b00000000 ;
			15'h000075F5 : data <= 8'b00000000 ;
			15'h000075F6 : data <= 8'b00000000 ;
			15'h000075F7 : data <= 8'b00000000 ;
			15'h000075F8 : data <= 8'b00000000 ;
			15'h000075F9 : data <= 8'b00000000 ;
			15'h000075FA : data <= 8'b00000000 ;
			15'h000075FB : data <= 8'b00000000 ;
			15'h000075FC : data <= 8'b00000000 ;
			15'h000075FD : data <= 8'b00000000 ;
			15'h000075FE : data <= 8'b00000000 ;
			15'h000075FF : data <= 8'b00000000 ;
			15'h00007600 : data <= 8'b00000000 ;
			15'h00007601 : data <= 8'b00000000 ;
			15'h00007602 : data <= 8'b00000000 ;
			15'h00007603 : data <= 8'b00000000 ;
			15'h00007604 : data <= 8'b00000000 ;
			15'h00007605 : data <= 8'b00000000 ;
			15'h00007606 : data <= 8'b00000000 ;
			15'h00007607 : data <= 8'b00000000 ;
			15'h00007608 : data <= 8'b00000000 ;
			15'h00007609 : data <= 8'b00000000 ;
			15'h0000760A : data <= 8'b00000000 ;
			15'h0000760B : data <= 8'b00000000 ;
			15'h0000760C : data <= 8'b00000000 ;
			15'h0000760D : data <= 8'b00000000 ;
			15'h0000760E : data <= 8'b00000000 ;
			15'h0000760F : data <= 8'b00000000 ;
			15'h00007610 : data <= 8'b00000000 ;
			15'h00007611 : data <= 8'b00000000 ;
			15'h00007612 : data <= 8'b00000000 ;
			15'h00007613 : data <= 8'b00000000 ;
			15'h00007614 : data <= 8'b00000000 ;
			15'h00007615 : data <= 8'b00000000 ;
			15'h00007616 : data <= 8'b00000000 ;
			15'h00007617 : data <= 8'b00000000 ;
			15'h00007618 : data <= 8'b00000000 ;
			15'h00007619 : data <= 8'b00000000 ;
			15'h0000761A : data <= 8'b00000000 ;
			15'h0000761B : data <= 8'b00000000 ;
			15'h0000761C : data <= 8'b00000000 ;
			15'h0000761D : data <= 8'b00000000 ;
			15'h0000761E : data <= 8'b00000000 ;
			15'h0000761F : data <= 8'b00000000 ;
			15'h00007620 : data <= 8'b00000000 ;
			15'h00007621 : data <= 8'b00000000 ;
			15'h00007622 : data <= 8'b00000000 ;
			15'h00007623 : data <= 8'b00000000 ;
			15'h00007624 : data <= 8'b00000000 ;
			15'h00007625 : data <= 8'b00000000 ;
			15'h00007626 : data <= 8'b00000000 ;
			15'h00007627 : data <= 8'b00000000 ;
			15'h00007628 : data <= 8'b00000000 ;
			15'h00007629 : data <= 8'b00000000 ;
			15'h0000762A : data <= 8'b00000000 ;
			15'h0000762B : data <= 8'b00000000 ;
			15'h0000762C : data <= 8'b00000000 ;
			15'h0000762D : data <= 8'b00000000 ;
			15'h0000762E : data <= 8'b00000000 ;
			15'h0000762F : data <= 8'b00000000 ;
			15'h00007630 : data <= 8'b00000000 ;
			15'h00007631 : data <= 8'b00000000 ;
			15'h00007632 : data <= 8'b00000000 ;
			15'h00007633 : data <= 8'b00000000 ;
			15'h00007634 : data <= 8'b00000000 ;
			15'h00007635 : data <= 8'b00000000 ;
			15'h00007636 : data <= 8'b00000000 ;
			15'h00007637 : data <= 8'b00000000 ;
			15'h00007638 : data <= 8'b00000000 ;
			15'h00007639 : data <= 8'b00000000 ;
			15'h0000763A : data <= 8'b00000000 ;
			15'h0000763B : data <= 8'b00000000 ;
			15'h0000763C : data <= 8'b00000000 ;
			15'h0000763D : data <= 8'b00000000 ;
			15'h0000763E : data <= 8'b00000000 ;
			15'h0000763F : data <= 8'b00000000 ;
			15'h00007640 : data <= 8'b00000000 ;
			15'h00007641 : data <= 8'b00000000 ;
			15'h00007642 : data <= 8'b00000000 ;
			15'h00007643 : data <= 8'b00000000 ;
			15'h00007644 : data <= 8'b00000000 ;
			15'h00007645 : data <= 8'b00000000 ;
			15'h00007646 : data <= 8'b00000000 ;
			15'h00007647 : data <= 8'b00000000 ;
			15'h00007648 : data <= 8'b00000000 ;
			15'h00007649 : data <= 8'b00000000 ;
			15'h0000764A : data <= 8'b00000000 ;
			15'h0000764B : data <= 8'b00000000 ;
			15'h0000764C : data <= 8'b00000000 ;
			15'h0000764D : data <= 8'b00000000 ;
			15'h0000764E : data <= 8'b00000000 ;
			15'h0000764F : data <= 8'b00000000 ;
			15'h00007650 : data <= 8'b00000000 ;
			15'h00007651 : data <= 8'b00000000 ;
			15'h00007652 : data <= 8'b00000000 ;
			15'h00007653 : data <= 8'b00000000 ;
			15'h00007654 : data <= 8'b00000000 ;
			15'h00007655 : data <= 8'b00000000 ;
			15'h00007656 : data <= 8'b00000000 ;
			15'h00007657 : data <= 8'b00000000 ;
			15'h00007658 : data <= 8'b00000000 ;
			15'h00007659 : data <= 8'b00000000 ;
			15'h0000765A : data <= 8'b00000000 ;
			15'h0000765B : data <= 8'b00000000 ;
			15'h0000765C : data <= 8'b00000000 ;
			15'h0000765D : data <= 8'b00000000 ;
			15'h0000765E : data <= 8'b00000000 ;
			15'h0000765F : data <= 8'b00000000 ;
			15'h00007660 : data <= 8'b00000000 ;
			15'h00007661 : data <= 8'b00000000 ;
			15'h00007662 : data <= 8'b00000000 ;
			15'h00007663 : data <= 8'b00000000 ;
			15'h00007664 : data <= 8'b00000000 ;
			15'h00007665 : data <= 8'b00000000 ;
			15'h00007666 : data <= 8'b00000000 ;
			15'h00007667 : data <= 8'b00000000 ;
			15'h00007668 : data <= 8'b00000000 ;
			15'h00007669 : data <= 8'b00000000 ;
			15'h0000766A : data <= 8'b00000000 ;
			15'h0000766B : data <= 8'b00000000 ;
			15'h0000766C : data <= 8'b00000000 ;
			15'h0000766D : data <= 8'b00000000 ;
			15'h0000766E : data <= 8'b00000000 ;
			15'h0000766F : data <= 8'b00000000 ;
			15'h00007670 : data <= 8'b00000000 ;
			15'h00007671 : data <= 8'b00000000 ;
			15'h00007672 : data <= 8'b00000000 ;
			15'h00007673 : data <= 8'b00000000 ;
			15'h00007674 : data <= 8'b00000000 ;
			15'h00007675 : data <= 8'b00000000 ;
			15'h00007676 : data <= 8'b00000000 ;
			15'h00007677 : data <= 8'b00000000 ;
			15'h00007678 : data <= 8'b00000000 ;
			15'h00007679 : data <= 8'b00000000 ;
			15'h0000767A : data <= 8'b00000000 ;
			15'h0000767B : data <= 8'b00000000 ;
			15'h0000767C : data <= 8'b00000000 ;
			15'h0000767D : data <= 8'b00000000 ;
			15'h0000767E : data <= 8'b00000000 ;
			15'h0000767F : data <= 8'b00000000 ;
			15'h00007680 : data <= 8'b00000000 ;
			15'h00007681 : data <= 8'b00000000 ;
			15'h00007682 : data <= 8'b00000000 ;
			15'h00007683 : data <= 8'b00000000 ;
			15'h00007684 : data <= 8'b00000000 ;
			15'h00007685 : data <= 8'b00000000 ;
			15'h00007686 : data <= 8'b00000000 ;
			15'h00007687 : data <= 8'b00000000 ;
			15'h00007688 : data <= 8'b00000000 ;
			15'h00007689 : data <= 8'b00000000 ;
			15'h0000768A : data <= 8'b00000000 ;
			15'h0000768B : data <= 8'b00000000 ;
			15'h0000768C : data <= 8'b00000000 ;
			15'h0000768D : data <= 8'b00000000 ;
			15'h0000768E : data <= 8'b00000000 ;
			15'h0000768F : data <= 8'b00000000 ;
			15'h00007690 : data <= 8'b00000000 ;
			15'h00007691 : data <= 8'b00000000 ;
			15'h00007692 : data <= 8'b00000000 ;
			15'h00007693 : data <= 8'b00000000 ;
			15'h00007694 : data <= 8'b00000000 ;
			15'h00007695 : data <= 8'b00000000 ;
			15'h00007696 : data <= 8'b00000000 ;
			15'h00007697 : data <= 8'b00000000 ;
			15'h00007698 : data <= 8'b00000000 ;
			15'h00007699 : data <= 8'b00000000 ;
			15'h0000769A : data <= 8'b00000000 ;
			15'h0000769B : data <= 8'b00000000 ;
			15'h0000769C : data <= 8'b00000000 ;
			15'h0000769D : data <= 8'b00000000 ;
			15'h0000769E : data <= 8'b00000000 ;
			15'h0000769F : data <= 8'b00000000 ;
			15'h000076A0 : data <= 8'b00000000 ;
			15'h000076A1 : data <= 8'b00000000 ;
			15'h000076A2 : data <= 8'b00000000 ;
			15'h000076A3 : data <= 8'b00000000 ;
			15'h000076A4 : data <= 8'b00000000 ;
			15'h000076A5 : data <= 8'b00000000 ;
			15'h000076A6 : data <= 8'b00000000 ;
			15'h000076A7 : data <= 8'b00000000 ;
			15'h000076A8 : data <= 8'b00000000 ;
			15'h000076A9 : data <= 8'b00000000 ;
			15'h000076AA : data <= 8'b00000000 ;
			15'h000076AB : data <= 8'b00000000 ;
			15'h000076AC : data <= 8'b00000000 ;
			15'h000076AD : data <= 8'b00000000 ;
			15'h000076AE : data <= 8'b00000000 ;
			15'h000076AF : data <= 8'b00000000 ;
			15'h000076B0 : data <= 8'b00000000 ;
			15'h000076B1 : data <= 8'b00000000 ;
			15'h000076B2 : data <= 8'b00000000 ;
			15'h000076B3 : data <= 8'b00000000 ;
			15'h000076B4 : data <= 8'b00000000 ;
			15'h000076B5 : data <= 8'b00000000 ;
			15'h000076B6 : data <= 8'b00000000 ;
			15'h000076B7 : data <= 8'b00000000 ;
			15'h000076B8 : data <= 8'b00000000 ;
			15'h000076B9 : data <= 8'b00000000 ;
			15'h000076BA : data <= 8'b00000000 ;
			15'h000076BB : data <= 8'b00000000 ;
			15'h000076BC : data <= 8'b00000000 ;
			15'h000076BD : data <= 8'b00000000 ;
			15'h000076BE : data <= 8'b00000000 ;
			15'h000076BF : data <= 8'b00000000 ;
			15'h000076C0 : data <= 8'b00000000 ;
			15'h000076C1 : data <= 8'b00000000 ;
			15'h000076C2 : data <= 8'b00000000 ;
			15'h000076C3 : data <= 8'b00000000 ;
			15'h000076C4 : data <= 8'b00000000 ;
			15'h000076C5 : data <= 8'b00000000 ;
			15'h000076C6 : data <= 8'b00000000 ;
			15'h000076C7 : data <= 8'b00000000 ;
			15'h000076C8 : data <= 8'b00000000 ;
			15'h000076C9 : data <= 8'b00000000 ;
			15'h000076CA : data <= 8'b00000000 ;
			15'h000076CB : data <= 8'b00000000 ;
			15'h000076CC : data <= 8'b00000000 ;
			15'h000076CD : data <= 8'b00000000 ;
			15'h000076CE : data <= 8'b00000000 ;
			15'h000076CF : data <= 8'b00000000 ;
			15'h000076D0 : data <= 8'b00000000 ;
			15'h000076D1 : data <= 8'b00000000 ;
			15'h000076D2 : data <= 8'b00000000 ;
			15'h000076D3 : data <= 8'b00000000 ;
			15'h000076D4 : data <= 8'b00000000 ;
			15'h000076D5 : data <= 8'b00000000 ;
			15'h000076D6 : data <= 8'b00000000 ;
			15'h000076D7 : data <= 8'b00000000 ;
			15'h000076D8 : data <= 8'b00000000 ;
			15'h000076D9 : data <= 8'b00000000 ;
			15'h000076DA : data <= 8'b00000000 ;
			15'h000076DB : data <= 8'b00000000 ;
			15'h000076DC : data <= 8'b00000000 ;
			15'h000076DD : data <= 8'b00000000 ;
			15'h000076DE : data <= 8'b00000000 ;
			15'h000076DF : data <= 8'b00000000 ;
			15'h000076E0 : data <= 8'b00000000 ;
			15'h000076E1 : data <= 8'b00000000 ;
			15'h000076E2 : data <= 8'b00000000 ;
			15'h000076E3 : data <= 8'b00000000 ;
			15'h000076E4 : data <= 8'b00000000 ;
			15'h000076E5 : data <= 8'b00000000 ;
			15'h000076E6 : data <= 8'b00000000 ;
			15'h000076E7 : data <= 8'b00000000 ;
			15'h000076E8 : data <= 8'b00000000 ;
			15'h000076E9 : data <= 8'b00000000 ;
			15'h000076EA : data <= 8'b00000000 ;
			15'h000076EB : data <= 8'b00000000 ;
			15'h000076EC : data <= 8'b00000000 ;
			15'h000076ED : data <= 8'b00000000 ;
			15'h000076EE : data <= 8'b00000000 ;
			15'h000076EF : data <= 8'b00000000 ;
			15'h000076F0 : data <= 8'b00000000 ;
			15'h000076F1 : data <= 8'b00000000 ;
			15'h000076F2 : data <= 8'b00000000 ;
			15'h000076F3 : data <= 8'b00000000 ;
			15'h000076F4 : data <= 8'b00000000 ;
			15'h000076F5 : data <= 8'b00000000 ;
			15'h000076F6 : data <= 8'b00000000 ;
			15'h000076F7 : data <= 8'b00000000 ;
			15'h000076F8 : data <= 8'b00000000 ;
			15'h000076F9 : data <= 8'b00000000 ;
			15'h000076FA : data <= 8'b00000000 ;
			15'h000076FB : data <= 8'b00000000 ;
			15'h000076FC : data <= 8'b00000000 ;
			15'h000076FD : data <= 8'b00000000 ;
			15'h000076FE : data <= 8'b00000000 ;
			15'h000076FF : data <= 8'b00000000 ;
			15'h00007700 : data <= 8'b00000000 ;
			15'h00007701 : data <= 8'b00000000 ;
			15'h00007702 : data <= 8'b00000000 ;
			15'h00007703 : data <= 8'b00000000 ;
			15'h00007704 : data <= 8'b00000000 ;
			15'h00007705 : data <= 8'b00000000 ;
			15'h00007706 : data <= 8'b00000000 ;
			15'h00007707 : data <= 8'b00000000 ;
			15'h00007708 : data <= 8'b00000000 ;
			15'h00007709 : data <= 8'b00000000 ;
			15'h0000770A : data <= 8'b00000000 ;
			15'h0000770B : data <= 8'b00000000 ;
			15'h0000770C : data <= 8'b00000000 ;
			15'h0000770D : data <= 8'b00000000 ;
			15'h0000770E : data <= 8'b00000000 ;
			15'h0000770F : data <= 8'b00000000 ;
			15'h00007710 : data <= 8'b00000000 ;
			15'h00007711 : data <= 8'b00000000 ;
			15'h00007712 : data <= 8'b00000000 ;
			15'h00007713 : data <= 8'b00000000 ;
			15'h00007714 : data <= 8'b00000000 ;
			15'h00007715 : data <= 8'b00000000 ;
			15'h00007716 : data <= 8'b00000000 ;
			15'h00007717 : data <= 8'b00000000 ;
			15'h00007718 : data <= 8'b00000000 ;
			15'h00007719 : data <= 8'b00000000 ;
			15'h0000771A : data <= 8'b00000000 ;
			15'h0000771B : data <= 8'b00000000 ;
			15'h0000771C : data <= 8'b00000000 ;
			15'h0000771D : data <= 8'b00000000 ;
			15'h0000771E : data <= 8'b00000000 ;
			15'h0000771F : data <= 8'b00000000 ;
			15'h00007720 : data <= 8'b00000000 ;
			15'h00007721 : data <= 8'b00000000 ;
			15'h00007722 : data <= 8'b00000000 ;
			15'h00007723 : data <= 8'b00000000 ;
			15'h00007724 : data <= 8'b00000000 ;
			15'h00007725 : data <= 8'b00000000 ;
			15'h00007726 : data <= 8'b00000000 ;
			15'h00007727 : data <= 8'b00000000 ;
			15'h00007728 : data <= 8'b00000000 ;
			15'h00007729 : data <= 8'b00000000 ;
			15'h0000772A : data <= 8'b00000000 ;
			15'h0000772B : data <= 8'b00000000 ;
			15'h0000772C : data <= 8'b00000000 ;
			15'h0000772D : data <= 8'b00000000 ;
			15'h0000772E : data <= 8'b00000000 ;
			15'h0000772F : data <= 8'b00000000 ;
			15'h00007730 : data <= 8'b00000000 ;
			15'h00007731 : data <= 8'b00000000 ;
			15'h00007732 : data <= 8'b00000000 ;
			15'h00007733 : data <= 8'b00000000 ;
			15'h00007734 : data <= 8'b00000000 ;
			15'h00007735 : data <= 8'b00000000 ;
			15'h00007736 : data <= 8'b00000000 ;
			15'h00007737 : data <= 8'b00000000 ;
			15'h00007738 : data <= 8'b00000000 ;
			15'h00007739 : data <= 8'b00000000 ;
			15'h0000773A : data <= 8'b00000000 ;
			15'h0000773B : data <= 8'b00000000 ;
			15'h0000773C : data <= 8'b00000000 ;
			15'h0000773D : data <= 8'b00000000 ;
			15'h0000773E : data <= 8'b00000000 ;
			15'h0000773F : data <= 8'b00000000 ;
			15'h00007740 : data <= 8'b00000000 ;
			15'h00007741 : data <= 8'b00000000 ;
			15'h00007742 : data <= 8'b00000000 ;
			15'h00007743 : data <= 8'b00000000 ;
			15'h00007744 : data <= 8'b00000000 ;
			15'h00007745 : data <= 8'b00000000 ;
			15'h00007746 : data <= 8'b00000000 ;
			15'h00007747 : data <= 8'b00000000 ;
			15'h00007748 : data <= 8'b00000000 ;
			15'h00007749 : data <= 8'b00000000 ;
			15'h0000774A : data <= 8'b00000000 ;
			15'h0000774B : data <= 8'b00000000 ;
			15'h0000774C : data <= 8'b00000000 ;
			15'h0000774D : data <= 8'b00000000 ;
			15'h0000774E : data <= 8'b00000000 ;
			15'h0000774F : data <= 8'b00000000 ;
			15'h00007750 : data <= 8'b00000000 ;
			15'h00007751 : data <= 8'b00000000 ;
			15'h00007752 : data <= 8'b00000000 ;
			15'h00007753 : data <= 8'b00000000 ;
			15'h00007754 : data <= 8'b00000000 ;
			15'h00007755 : data <= 8'b00000000 ;
			15'h00007756 : data <= 8'b00000000 ;
			15'h00007757 : data <= 8'b00000000 ;
			15'h00007758 : data <= 8'b00000000 ;
			15'h00007759 : data <= 8'b00000000 ;
			15'h0000775A : data <= 8'b00000000 ;
			15'h0000775B : data <= 8'b00000000 ;
			15'h0000775C : data <= 8'b00000000 ;
			15'h0000775D : data <= 8'b00000000 ;
			15'h0000775E : data <= 8'b00000000 ;
			15'h0000775F : data <= 8'b00000000 ;
			15'h00007760 : data <= 8'b00000000 ;
			15'h00007761 : data <= 8'b00000000 ;
			15'h00007762 : data <= 8'b00000000 ;
			15'h00007763 : data <= 8'b00000000 ;
			15'h00007764 : data <= 8'b00000000 ;
			15'h00007765 : data <= 8'b00000000 ;
			15'h00007766 : data <= 8'b00000000 ;
			15'h00007767 : data <= 8'b00000000 ;
			15'h00007768 : data <= 8'b00000000 ;
			15'h00007769 : data <= 8'b00000000 ;
			15'h0000776A : data <= 8'b00000000 ;
			15'h0000776B : data <= 8'b00000000 ;
			15'h0000776C : data <= 8'b00000000 ;
			15'h0000776D : data <= 8'b00000000 ;
			15'h0000776E : data <= 8'b00000000 ;
			15'h0000776F : data <= 8'b00000000 ;
			15'h00007770 : data <= 8'b00000000 ;
			15'h00007771 : data <= 8'b00000000 ;
			15'h00007772 : data <= 8'b00000000 ;
			15'h00007773 : data <= 8'b00000000 ;
			15'h00007774 : data <= 8'b00000000 ;
			15'h00007775 : data <= 8'b00000000 ;
			15'h00007776 : data <= 8'b00000000 ;
			15'h00007777 : data <= 8'b00000000 ;
			15'h00007778 : data <= 8'b00000000 ;
			15'h00007779 : data <= 8'b00000000 ;
			15'h0000777A : data <= 8'b00000000 ;
			15'h0000777B : data <= 8'b00000000 ;
			15'h0000777C : data <= 8'b00000000 ;
			15'h0000777D : data <= 8'b00000000 ;
			15'h0000777E : data <= 8'b00000000 ;
			15'h0000777F : data <= 8'b00000000 ;
			15'h00007780 : data <= 8'b00000000 ;
			15'h00007781 : data <= 8'b00000000 ;
			15'h00007782 : data <= 8'b00000000 ;
			15'h00007783 : data <= 8'b00000000 ;
			15'h00007784 : data <= 8'b00000000 ;
			15'h00007785 : data <= 8'b00000000 ;
			15'h00007786 : data <= 8'b00000000 ;
			15'h00007787 : data <= 8'b00000000 ;
			15'h00007788 : data <= 8'b00000000 ;
			15'h00007789 : data <= 8'b00000000 ;
			15'h0000778A : data <= 8'b00000000 ;
			15'h0000778B : data <= 8'b00000000 ;
			15'h0000778C : data <= 8'b00000000 ;
			15'h0000778D : data <= 8'b00000000 ;
			15'h0000778E : data <= 8'b00000000 ;
			15'h0000778F : data <= 8'b00000000 ;
			15'h00007790 : data <= 8'b00000000 ;
			15'h00007791 : data <= 8'b00000000 ;
			15'h00007792 : data <= 8'b00000000 ;
			15'h00007793 : data <= 8'b00000000 ;
			15'h00007794 : data <= 8'b00000000 ;
			15'h00007795 : data <= 8'b00000000 ;
			15'h00007796 : data <= 8'b00000000 ;
			15'h00007797 : data <= 8'b00000000 ;
			15'h00007798 : data <= 8'b00000000 ;
			15'h00007799 : data <= 8'b00000000 ;
			15'h0000779A : data <= 8'b00000000 ;
			15'h0000779B : data <= 8'b00000000 ;
			15'h0000779C : data <= 8'b00000000 ;
			15'h0000779D : data <= 8'b00000000 ;
			15'h0000779E : data <= 8'b00000000 ;
			15'h0000779F : data <= 8'b00000000 ;
			15'h000077A0 : data <= 8'b00000000 ;
			15'h000077A1 : data <= 8'b00000000 ;
			15'h000077A2 : data <= 8'b00000000 ;
			15'h000077A3 : data <= 8'b00000000 ;
			15'h000077A4 : data <= 8'b00000000 ;
			15'h000077A5 : data <= 8'b00000000 ;
			15'h000077A6 : data <= 8'b00000000 ;
			15'h000077A7 : data <= 8'b00000000 ;
			15'h000077A8 : data <= 8'b00000000 ;
			15'h000077A9 : data <= 8'b00000000 ;
			15'h000077AA : data <= 8'b00000000 ;
			15'h000077AB : data <= 8'b00000000 ;
			15'h000077AC : data <= 8'b00000000 ;
			15'h000077AD : data <= 8'b00000000 ;
			15'h000077AE : data <= 8'b00000000 ;
			15'h000077AF : data <= 8'b00000000 ;
			15'h000077B0 : data <= 8'b00000000 ;
			15'h000077B1 : data <= 8'b00000000 ;
			15'h000077B2 : data <= 8'b00000000 ;
			15'h000077B3 : data <= 8'b00000000 ;
			15'h000077B4 : data <= 8'b00000000 ;
			15'h000077B5 : data <= 8'b00000000 ;
			15'h000077B6 : data <= 8'b00000000 ;
			15'h000077B7 : data <= 8'b00000000 ;
			15'h000077B8 : data <= 8'b00000000 ;
			15'h000077B9 : data <= 8'b00000000 ;
			15'h000077BA : data <= 8'b00000000 ;
			15'h000077BB : data <= 8'b00000000 ;
			15'h000077BC : data <= 8'b00000000 ;
			15'h000077BD : data <= 8'b00000000 ;
			15'h000077BE : data <= 8'b00000000 ;
			15'h000077BF : data <= 8'b00000000 ;
			15'h000077C0 : data <= 8'b00000000 ;
			15'h000077C1 : data <= 8'b00000000 ;
			15'h000077C2 : data <= 8'b00000000 ;
			15'h000077C3 : data <= 8'b00000000 ;
			15'h000077C4 : data <= 8'b00000000 ;
			15'h000077C5 : data <= 8'b00000000 ;
			15'h000077C6 : data <= 8'b00000000 ;
			15'h000077C7 : data <= 8'b00000000 ;
			15'h000077C8 : data <= 8'b00000000 ;
			15'h000077C9 : data <= 8'b00000000 ;
			15'h000077CA : data <= 8'b00000000 ;
			15'h000077CB : data <= 8'b00000000 ;
			15'h000077CC : data <= 8'b00000000 ;
			15'h000077CD : data <= 8'b00000000 ;
			15'h000077CE : data <= 8'b00000000 ;
			15'h000077CF : data <= 8'b00000000 ;
			15'h000077D0 : data <= 8'b00000000 ;
			15'h000077D1 : data <= 8'b00000000 ;
			15'h000077D2 : data <= 8'b00000000 ;
			15'h000077D3 : data <= 8'b00000000 ;
			15'h000077D4 : data <= 8'b00000000 ;
			15'h000077D5 : data <= 8'b00000000 ;
			15'h000077D6 : data <= 8'b00000000 ;
			15'h000077D7 : data <= 8'b00000000 ;
			15'h000077D8 : data <= 8'b00000000 ;
			15'h000077D9 : data <= 8'b00000000 ;
			15'h000077DA : data <= 8'b00000000 ;
			15'h000077DB : data <= 8'b00000000 ;
			15'h000077DC : data <= 8'b00000000 ;
			15'h000077DD : data <= 8'b00000000 ;
			15'h000077DE : data <= 8'b00000000 ;
			15'h000077DF : data <= 8'b00000000 ;
			15'h000077E0 : data <= 8'b00000000 ;
			15'h000077E1 : data <= 8'b00000000 ;
			15'h000077E2 : data <= 8'b00000000 ;
			15'h000077E3 : data <= 8'b00000000 ;
			15'h000077E4 : data <= 8'b00000000 ;
			15'h000077E5 : data <= 8'b00000000 ;
			15'h000077E6 : data <= 8'b00000000 ;
			15'h000077E7 : data <= 8'b00000000 ;
			15'h000077E8 : data <= 8'b00000000 ;
			15'h000077E9 : data <= 8'b00000000 ;
			15'h000077EA : data <= 8'b00000000 ;
			15'h000077EB : data <= 8'b00000000 ;
			15'h000077EC : data <= 8'b00000000 ;
			15'h000077ED : data <= 8'b00000000 ;
			15'h000077EE : data <= 8'b00000000 ;
			15'h000077EF : data <= 8'b00000000 ;
			15'h000077F0 : data <= 8'b00000000 ;
			15'h000077F1 : data <= 8'b00000000 ;
			15'h000077F2 : data <= 8'b00000000 ;
			15'h000077F3 : data <= 8'b00000000 ;
			15'h000077F4 : data <= 8'b00000000 ;
			15'h000077F5 : data <= 8'b00000000 ;
			15'h000077F6 : data <= 8'b00000000 ;
			15'h000077F7 : data <= 8'b00000000 ;
			15'h000077F8 : data <= 8'b00000000 ;
			15'h000077F9 : data <= 8'b00000000 ;
			15'h000077FA : data <= 8'b00000000 ;
			15'h000077FB : data <= 8'b00000000 ;
			15'h000077FC : data <= 8'b00000000 ;
			15'h000077FD : data <= 8'b00000000 ;
			15'h000077FE : data <= 8'b00000000 ;
			15'h000077FF : data <= 8'b00000000 ;
			15'h00007800 : data <= 8'b00000000 ;
			15'h00007801 : data <= 8'b00000000 ;
			15'h00007802 : data <= 8'b00000000 ;
			15'h00007803 : data <= 8'b00000000 ;
			15'h00007804 : data <= 8'b00000000 ;
			15'h00007805 : data <= 8'b00000000 ;
			15'h00007806 : data <= 8'b00000000 ;
			15'h00007807 : data <= 8'b00000000 ;
			15'h00007808 : data <= 8'b00000000 ;
			15'h00007809 : data <= 8'b00000000 ;
			15'h0000780A : data <= 8'b00000000 ;
			15'h0000780B : data <= 8'b00000000 ;
			15'h0000780C : data <= 8'b00000000 ;
			15'h0000780D : data <= 8'b00000000 ;
			15'h0000780E : data <= 8'b00000000 ;
			15'h0000780F : data <= 8'b00000000 ;
			15'h00007810 : data <= 8'b00000000 ;
			15'h00007811 : data <= 8'b00000000 ;
			15'h00007812 : data <= 8'b00000000 ;
			15'h00007813 : data <= 8'b00000000 ;
			15'h00007814 : data <= 8'b00000000 ;
			15'h00007815 : data <= 8'b00000000 ;
			15'h00007816 : data <= 8'b00000000 ;
			15'h00007817 : data <= 8'b00000000 ;
			15'h00007818 : data <= 8'b00000000 ;
			15'h00007819 : data <= 8'b00000000 ;
			15'h0000781A : data <= 8'b00000000 ;
			15'h0000781B : data <= 8'b00000000 ;
			15'h0000781C : data <= 8'b00000000 ;
			15'h0000781D : data <= 8'b00000000 ;
			15'h0000781E : data <= 8'b00000000 ;
			15'h0000781F : data <= 8'b00000000 ;
			15'h00007820 : data <= 8'b00000000 ;
			15'h00007821 : data <= 8'b00000000 ;
			15'h00007822 : data <= 8'b00000000 ;
			15'h00007823 : data <= 8'b00000000 ;
			15'h00007824 : data <= 8'b00000000 ;
			15'h00007825 : data <= 8'b00000000 ;
			15'h00007826 : data <= 8'b00000000 ;
			15'h00007827 : data <= 8'b00000000 ;
			15'h00007828 : data <= 8'b00000000 ;
			15'h00007829 : data <= 8'b00000000 ;
			15'h0000782A : data <= 8'b00000000 ;
			15'h0000782B : data <= 8'b00000000 ;
			15'h0000782C : data <= 8'b00000000 ;
			15'h0000782D : data <= 8'b00000000 ;
			15'h0000782E : data <= 8'b00000000 ;
			15'h0000782F : data <= 8'b00000000 ;
			15'h00007830 : data <= 8'b00000000 ;
			15'h00007831 : data <= 8'b00000000 ;
			15'h00007832 : data <= 8'b00000000 ;
			15'h00007833 : data <= 8'b00000000 ;
			15'h00007834 : data <= 8'b00000000 ;
			15'h00007835 : data <= 8'b00000000 ;
			15'h00007836 : data <= 8'b00000000 ;
			15'h00007837 : data <= 8'b00000000 ;
			15'h00007838 : data <= 8'b00000000 ;
			15'h00007839 : data <= 8'b00000000 ;
			15'h0000783A : data <= 8'b00000000 ;
			15'h0000783B : data <= 8'b00000000 ;
			15'h0000783C : data <= 8'b00000000 ;
			15'h0000783D : data <= 8'b00000000 ;
			15'h0000783E : data <= 8'b00000000 ;
			15'h0000783F : data <= 8'b00000000 ;
			15'h00007840 : data <= 8'b00000000 ;
			15'h00007841 : data <= 8'b00000000 ;
			15'h00007842 : data <= 8'b00000000 ;
			15'h00007843 : data <= 8'b00000000 ;
			15'h00007844 : data <= 8'b00000000 ;
			15'h00007845 : data <= 8'b00000000 ;
			15'h00007846 : data <= 8'b00000000 ;
			15'h00007847 : data <= 8'b00000000 ;
			15'h00007848 : data <= 8'b00000000 ;
			15'h00007849 : data <= 8'b00000000 ;
			15'h0000784A : data <= 8'b00000000 ;
			15'h0000784B : data <= 8'b00000000 ;
			15'h0000784C : data <= 8'b00000000 ;
			15'h0000784D : data <= 8'b00000000 ;
			15'h0000784E : data <= 8'b00000000 ;
			15'h0000784F : data <= 8'b00000000 ;
			15'h00007850 : data <= 8'b00000000 ;
			15'h00007851 : data <= 8'b00000000 ;
			15'h00007852 : data <= 8'b00000000 ;
			15'h00007853 : data <= 8'b00000000 ;
			15'h00007854 : data <= 8'b00000000 ;
			15'h00007855 : data <= 8'b00000000 ;
			15'h00007856 : data <= 8'b00000000 ;
			15'h00007857 : data <= 8'b00000000 ;
			15'h00007858 : data <= 8'b00000000 ;
			15'h00007859 : data <= 8'b00000000 ;
			15'h0000785A : data <= 8'b00000000 ;
			15'h0000785B : data <= 8'b00000000 ;
			15'h0000785C : data <= 8'b00000000 ;
			15'h0000785D : data <= 8'b00000000 ;
			15'h0000785E : data <= 8'b00000000 ;
			15'h0000785F : data <= 8'b00000000 ;
			15'h00007860 : data <= 8'b00000000 ;
			15'h00007861 : data <= 8'b00000000 ;
			15'h00007862 : data <= 8'b00000000 ;
			15'h00007863 : data <= 8'b00000000 ;
			15'h00007864 : data <= 8'b00000000 ;
			15'h00007865 : data <= 8'b00000000 ;
			15'h00007866 : data <= 8'b00000000 ;
			15'h00007867 : data <= 8'b00000000 ;
			15'h00007868 : data <= 8'b00000000 ;
			15'h00007869 : data <= 8'b00000000 ;
			15'h0000786A : data <= 8'b00000000 ;
			15'h0000786B : data <= 8'b00000000 ;
			15'h0000786C : data <= 8'b00000000 ;
			15'h0000786D : data <= 8'b00000000 ;
			15'h0000786E : data <= 8'b00000000 ;
			15'h0000786F : data <= 8'b00000000 ;
			15'h00007870 : data <= 8'b00000000 ;
			15'h00007871 : data <= 8'b00000000 ;
			15'h00007872 : data <= 8'b00000000 ;
			15'h00007873 : data <= 8'b00000000 ;
			15'h00007874 : data <= 8'b00000000 ;
			15'h00007875 : data <= 8'b00000000 ;
			15'h00007876 : data <= 8'b00000000 ;
			15'h00007877 : data <= 8'b00000000 ;
			15'h00007878 : data <= 8'b00000000 ;
			15'h00007879 : data <= 8'b00000000 ;
			15'h0000787A : data <= 8'b00000000 ;
			15'h0000787B : data <= 8'b00000000 ;
			15'h0000787C : data <= 8'b00000000 ;
			15'h0000787D : data <= 8'b00000000 ;
			15'h0000787E : data <= 8'b00000000 ;
			15'h0000787F : data <= 8'b00000000 ;
			15'h00007880 : data <= 8'b00000000 ;
			15'h00007881 : data <= 8'b00000000 ;
			15'h00007882 : data <= 8'b00000000 ;
			15'h00007883 : data <= 8'b00000000 ;
			15'h00007884 : data <= 8'b00000000 ;
			15'h00007885 : data <= 8'b00000000 ;
			15'h00007886 : data <= 8'b00000000 ;
			15'h00007887 : data <= 8'b00000000 ;
			15'h00007888 : data <= 8'b00000000 ;
			15'h00007889 : data <= 8'b00000000 ;
			15'h0000788A : data <= 8'b00000000 ;
			15'h0000788B : data <= 8'b00000000 ;
			15'h0000788C : data <= 8'b00000000 ;
			15'h0000788D : data <= 8'b00000000 ;
			15'h0000788E : data <= 8'b00000000 ;
			15'h0000788F : data <= 8'b00000000 ;
			15'h00007890 : data <= 8'b00000000 ;
			15'h00007891 : data <= 8'b00000000 ;
			15'h00007892 : data <= 8'b00000000 ;
			15'h00007893 : data <= 8'b00000000 ;
			15'h00007894 : data <= 8'b00000000 ;
			15'h00007895 : data <= 8'b00000000 ;
			15'h00007896 : data <= 8'b00000000 ;
			15'h00007897 : data <= 8'b00000000 ;
			15'h00007898 : data <= 8'b00000000 ;
			15'h00007899 : data <= 8'b00000000 ;
			15'h0000789A : data <= 8'b00000000 ;
			15'h0000789B : data <= 8'b00000000 ;
			15'h0000789C : data <= 8'b00000000 ;
			15'h0000789D : data <= 8'b00000000 ;
			15'h0000789E : data <= 8'b00000000 ;
			15'h0000789F : data <= 8'b00000000 ;
			15'h000078A0 : data <= 8'b00000000 ;
			15'h000078A1 : data <= 8'b00000000 ;
			15'h000078A2 : data <= 8'b00000000 ;
			15'h000078A3 : data <= 8'b00000000 ;
			15'h000078A4 : data <= 8'b00000000 ;
			15'h000078A5 : data <= 8'b00000000 ;
			15'h000078A6 : data <= 8'b00000000 ;
			15'h000078A7 : data <= 8'b00000000 ;
			15'h000078A8 : data <= 8'b00000000 ;
			15'h000078A9 : data <= 8'b00000000 ;
			15'h000078AA : data <= 8'b00000000 ;
			15'h000078AB : data <= 8'b00000000 ;
			15'h000078AC : data <= 8'b00000000 ;
			15'h000078AD : data <= 8'b00000000 ;
			15'h000078AE : data <= 8'b00000000 ;
			15'h000078AF : data <= 8'b00000000 ;
			15'h000078B0 : data <= 8'b00000000 ;
			15'h000078B1 : data <= 8'b00000000 ;
			15'h000078B2 : data <= 8'b00000000 ;
			15'h000078B3 : data <= 8'b00000000 ;
			15'h000078B4 : data <= 8'b00000000 ;
			15'h000078B5 : data <= 8'b00000000 ;
			15'h000078B6 : data <= 8'b00000000 ;
			15'h000078B7 : data <= 8'b00000000 ;
			15'h000078B8 : data <= 8'b00000000 ;
			15'h000078B9 : data <= 8'b00000000 ;
			15'h000078BA : data <= 8'b00000000 ;
			15'h000078BB : data <= 8'b00000000 ;
			15'h000078BC : data <= 8'b00000000 ;
			15'h000078BD : data <= 8'b00000000 ;
			15'h000078BE : data <= 8'b00000000 ;
			15'h000078BF : data <= 8'b00000000 ;
			15'h000078C0 : data <= 8'b00000000 ;
			15'h000078C1 : data <= 8'b00000000 ;
			15'h000078C2 : data <= 8'b00000000 ;
			15'h000078C3 : data <= 8'b00000000 ;
			15'h000078C4 : data <= 8'b00000000 ;
			15'h000078C5 : data <= 8'b00000000 ;
			15'h000078C6 : data <= 8'b00000000 ;
			15'h000078C7 : data <= 8'b00000000 ;
			15'h000078C8 : data <= 8'b00000000 ;
			15'h000078C9 : data <= 8'b00000000 ;
			15'h000078CA : data <= 8'b00000000 ;
			15'h000078CB : data <= 8'b00000000 ;
			15'h000078CC : data <= 8'b00000000 ;
			15'h000078CD : data <= 8'b00000000 ;
			15'h000078CE : data <= 8'b00000000 ;
			15'h000078CF : data <= 8'b00000000 ;
			15'h000078D0 : data <= 8'b00000000 ;
			15'h000078D1 : data <= 8'b00000000 ;
			15'h000078D2 : data <= 8'b00000000 ;
			15'h000078D3 : data <= 8'b00000000 ;
			15'h000078D4 : data <= 8'b00000000 ;
			15'h000078D5 : data <= 8'b00000000 ;
			15'h000078D6 : data <= 8'b00000000 ;
			15'h000078D7 : data <= 8'b00000000 ;
			15'h000078D8 : data <= 8'b00000000 ;
			15'h000078D9 : data <= 8'b00000000 ;
			15'h000078DA : data <= 8'b00000000 ;
			15'h000078DB : data <= 8'b00000000 ;
			15'h000078DC : data <= 8'b00000000 ;
			15'h000078DD : data <= 8'b00000000 ;
			15'h000078DE : data <= 8'b00000000 ;
			15'h000078DF : data <= 8'b00000000 ;
			15'h000078E0 : data <= 8'b00000000 ;
			15'h000078E1 : data <= 8'b00000000 ;
			15'h000078E2 : data <= 8'b00000000 ;
			15'h000078E3 : data <= 8'b00000000 ;
			15'h000078E4 : data <= 8'b00000000 ;
			15'h000078E5 : data <= 8'b00000000 ;
			15'h000078E6 : data <= 8'b00000000 ;
			15'h000078E7 : data <= 8'b00000000 ;
			15'h000078E8 : data <= 8'b00000000 ;
			15'h000078E9 : data <= 8'b00000000 ;
			15'h000078EA : data <= 8'b00000000 ;
			15'h000078EB : data <= 8'b00000000 ;
			15'h000078EC : data <= 8'b00000000 ;
			15'h000078ED : data <= 8'b00000000 ;
			15'h000078EE : data <= 8'b00000000 ;
			15'h000078EF : data <= 8'b00000000 ;
			15'h000078F0 : data <= 8'b00000000 ;
			15'h000078F1 : data <= 8'b00000000 ;
			15'h000078F2 : data <= 8'b00000000 ;
			15'h000078F3 : data <= 8'b00000000 ;
			15'h000078F4 : data <= 8'b00000000 ;
			15'h000078F5 : data <= 8'b00000000 ;
			15'h000078F6 : data <= 8'b00000000 ;
			15'h000078F7 : data <= 8'b00000000 ;
			15'h000078F8 : data <= 8'b00000000 ;
			15'h000078F9 : data <= 8'b00000000 ;
			15'h000078FA : data <= 8'b00000000 ;
			15'h000078FB : data <= 8'b00000000 ;
			15'h000078FC : data <= 8'b00000000 ;
			15'h000078FD : data <= 8'b00000000 ;
			15'h000078FE : data <= 8'b00000000 ;
			15'h000078FF : data <= 8'b00000000 ;
			15'h00007900 : data <= 8'b00000000 ;
			15'h00007901 : data <= 8'b00000000 ;
			15'h00007902 : data <= 8'b00000000 ;
			15'h00007903 : data <= 8'b00000000 ;
			15'h00007904 : data <= 8'b00000000 ;
			15'h00007905 : data <= 8'b00000000 ;
			15'h00007906 : data <= 8'b00000000 ;
			15'h00007907 : data <= 8'b00000000 ;
			15'h00007908 : data <= 8'b00000000 ;
			15'h00007909 : data <= 8'b00000000 ;
			15'h0000790A : data <= 8'b00000000 ;
			15'h0000790B : data <= 8'b00000000 ;
			15'h0000790C : data <= 8'b00000000 ;
			15'h0000790D : data <= 8'b00000000 ;
			15'h0000790E : data <= 8'b00000000 ;
			15'h0000790F : data <= 8'b00000000 ;
			15'h00007910 : data <= 8'b00000000 ;
			15'h00007911 : data <= 8'b00000000 ;
			15'h00007912 : data <= 8'b00000000 ;
			15'h00007913 : data <= 8'b00000000 ;
			15'h00007914 : data <= 8'b00000000 ;
			15'h00007915 : data <= 8'b00000000 ;
			15'h00007916 : data <= 8'b00000000 ;
			15'h00007917 : data <= 8'b00000000 ;
			15'h00007918 : data <= 8'b00000000 ;
			15'h00007919 : data <= 8'b00000000 ;
			15'h0000791A : data <= 8'b00000000 ;
			15'h0000791B : data <= 8'b00000000 ;
			15'h0000791C : data <= 8'b00000000 ;
			15'h0000791D : data <= 8'b00000000 ;
			15'h0000791E : data <= 8'b00000000 ;
			15'h0000791F : data <= 8'b00000000 ;
			15'h00007920 : data <= 8'b00000000 ;
			15'h00007921 : data <= 8'b00000000 ;
			15'h00007922 : data <= 8'b00000000 ;
			15'h00007923 : data <= 8'b00000000 ;
			15'h00007924 : data <= 8'b00000000 ;
			15'h00007925 : data <= 8'b00000000 ;
			15'h00007926 : data <= 8'b00000000 ;
			15'h00007927 : data <= 8'b00000000 ;
			15'h00007928 : data <= 8'b00000000 ;
			15'h00007929 : data <= 8'b00000000 ;
			15'h0000792A : data <= 8'b00000000 ;
			15'h0000792B : data <= 8'b00000000 ;
			15'h0000792C : data <= 8'b00000000 ;
			15'h0000792D : data <= 8'b00000000 ;
			15'h0000792E : data <= 8'b00000000 ;
			15'h0000792F : data <= 8'b00000000 ;
			15'h00007930 : data <= 8'b00000000 ;
			15'h00007931 : data <= 8'b00000000 ;
			15'h00007932 : data <= 8'b00000000 ;
			15'h00007933 : data <= 8'b00000000 ;
			15'h00007934 : data <= 8'b00000000 ;
			15'h00007935 : data <= 8'b00000000 ;
			15'h00007936 : data <= 8'b00000000 ;
			15'h00007937 : data <= 8'b00000000 ;
			15'h00007938 : data <= 8'b00000000 ;
			15'h00007939 : data <= 8'b00000000 ;
			15'h0000793A : data <= 8'b00000000 ;
			15'h0000793B : data <= 8'b00000000 ;
			15'h0000793C : data <= 8'b00000000 ;
			15'h0000793D : data <= 8'b00000000 ;
			15'h0000793E : data <= 8'b00000000 ;
			15'h0000793F : data <= 8'b00000000 ;
			15'h00007940 : data <= 8'b00000000 ;
			15'h00007941 : data <= 8'b00000000 ;
			15'h00007942 : data <= 8'b00000000 ;
			15'h00007943 : data <= 8'b00000000 ;
			15'h00007944 : data <= 8'b00000000 ;
			15'h00007945 : data <= 8'b00000000 ;
			15'h00007946 : data <= 8'b00000000 ;
			15'h00007947 : data <= 8'b00000000 ;
			15'h00007948 : data <= 8'b00000000 ;
			15'h00007949 : data <= 8'b00000000 ;
			15'h0000794A : data <= 8'b00000000 ;
			15'h0000794B : data <= 8'b00000000 ;
			15'h0000794C : data <= 8'b00000000 ;
			15'h0000794D : data <= 8'b00000000 ;
			15'h0000794E : data <= 8'b00000000 ;
			15'h0000794F : data <= 8'b00000000 ;
			15'h00007950 : data <= 8'b00000000 ;
			15'h00007951 : data <= 8'b00000000 ;
			15'h00007952 : data <= 8'b00000000 ;
			15'h00007953 : data <= 8'b00000000 ;
			15'h00007954 : data <= 8'b00000000 ;
			15'h00007955 : data <= 8'b00000000 ;
			15'h00007956 : data <= 8'b00000000 ;
			15'h00007957 : data <= 8'b00000000 ;
			15'h00007958 : data <= 8'b00000000 ;
			15'h00007959 : data <= 8'b00000000 ;
			15'h0000795A : data <= 8'b00000000 ;
			15'h0000795B : data <= 8'b00000000 ;
			15'h0000795C : data <= 8'b00000000 ;
			15'h0000795D : data <= 8'b00000000 ;
			15'h0000795E : data <= 8'b00000000 ;
			15'h0000795F : data <= 8'b00000000 ;
			15'h00007960 : data <= 8'b00000000 ;
			15'h00007961 : data <= 8'b00000000 ;
			15'h00007962 : data <= 8'b00000000 ;
			15'h00007963 : data <= 8'b00000000 ;
			15'h00007964 : data <= 8'b00000000 ;
			15'h00007965 : data <= 8'b00000000 ;
			15'h00007966 : data <= 8'b00000000 ;
			15'h00007967 : data <= 8'b00000000 ;
			15'h00007968 : data <= 8'b00000000 ;
			15'h00007969 : data <= 8'b00000000 ;
			15'h0000796A : data <= 8'b00000000 ;
			15'h0000796B : data <= 8'b00000000 ;
			15'h0000796C : data <= 8'b00000000 ;
			15'h0000796D : data <= 8'b00000000 ;
			15'h0000796E : data <= 8'b00000000 ;
			15'h0000796F : data <= 8'b00000000 ;
			15'h00007970 : data <= 8'b00000000 ;
			15'h00007971 : data <= 8'b00000000 ;
			15'h00007972 : data <= 8'b00000000 ;
			15'h00007973 : data <= 8'b00000000 ;
			15'h00007974 : data <= 8'b00000000 ;
			15'h00007975 : data <= 8'b00000000 ;
			15'h00007976 : data <= 8'b00000000 ;
			15'h00007977 : data <= 8'b00000000 ;
			15'h00007978 : data <= 8'b00000000 ;
			15'h00007979 : data <= 8'b00000000 ;
			15'h0000797A : data <= 8'b00000000 ;
			15'h0000797B : data <= 8'b00000000 ;
			15'h0000797C : data <= 8'b00000000 ;
			15'h0000797D : data <= 8'b00000000 ;
			15'h0000797E : data <= 8'b00000000 ;
			15'h0000797F : data <= 8'b00000000 ;
			15'h00007980 : data <= 8'b00000000 ;
			15'h00007981 : data <= 8'b00000000 ;
			15'h00007982 : data <= 8'b00000000 ;
			15'h00007983 : data <= 8'b00000000 ;
			15'h00007984 : data <= 8'b00000000 ;
			15'h00007985 : data <= 8'b00000000 ;
			15'h00007986 : data <= 8'b00000000 ;
			15'h00007987 : data <= 8'b00000000 ;
			15'h00007988 : data <= 8'b00000000 ;
			15'h00007989 : data <= 8'b00000000 ;
			15'h0000798A : data <= 8'b00000000 ;
			15'h0000798B : data <= 8'b00000000 ;
			15'h0000798C : data <= 8'b00000000 ;
			15'h0000798D : data <= 8'b00000000 ;
			15'h0000798E : data <= 8'b00000000 ;
			15'h0000798F : data <= 8'b00000000 ;
			15'h00007990 : data <= 8'b00000000 ;
			15'h00007991 : data <= 8'b00000000 ;
			15'h00007992 : data <= 8'b00000000 ;
			15'h00007993 : data <= 8'b00000000 ;
			15'h00007994 : data <= 8'b00000000 ;
			15'h00007995 : data <= 8'b00000000 ;
			15'h00007996 : data <= 8'b00000000 ;
			15'h00007997 : data <= 8'b00000000 ;
			15'h00007998 : data <= 8'b00000000 ;
			15'h00007999 : data <= 8'b00000000 ;
			15'h0000799A : data <= 8'b00000000 ;
			15'h0000799B : data <= 8'b00000000 ;
			15'h0000799C : data <= 8'b00000000 ;
			15'h0000799D : data <= 8'b00000000 ;
			15'h0000799E : data <= 8'b00000000 ;
			15'h0000799F : data <= 8'b00000000 ;
			15'h000079A0 : data <= 8'b00000000 ;
			15'h000079A1 : data <= 8'b00000000 ;
			15'h000079A2 : data <= 8'b00000000 ;
			15'h000079A3 : data <= 8'b00000000 ;
			15'h000079A4 : data <= 8'b00000000 ;
			15'h000079A5 : data <= 8'b00000000 ;
			15'h000079A6 : data <= 8'b00000000 ;
			15'h000079A7 : data <= 8'b00000000 ;
			15'h000079A8 : data <= 8'b00000000 ;
			15'h000079A9 : data <= 8'b00000000 ;
			15'h000079AA : data <= 8'b00000000 ;
			15'h000079AB : data <= 8'b00000000 ;
			15'h000079AC : data <= 8'b00000000 ;
			15'h000079AD : data <= 8'b00000000 ;
			15'h000079AE : data <= 8'b00000000 ;
			15'h000079AF : data <= 8'b00000000 ;
			15'h000079B0 : data <= 8'b00000000 ;
			15'h000079B1 : data <= 8'b00000000 ;
			15'h000079B2 : data <= 8'b00000000 ;
			15'h000079B3 : data <= 8'b00000000 ;
			15'h000079B4 : data <= 8'b00000000 ;
			15'h000079B5 : data <= 8'b00000000 ;
			15'h000079B6 : data <= 8'b00000000 ;
			15'h000079B7 : data <= 8'b00000000 ;
			15'h000079B8 : data <= 8'b00000000 ;
			15'h000079B9 : data <= 8'b00000000 ;
			15'h000079BA : data <= 8'b00000000 ;
			15'h000079BB : data <= 8'b00000000 ;
			15'h000079BC : data <= 8'b00000000 ;
			15'h000079BD : data <= 8'b00000000 ;
			15'h000079BE : data <= 8'b00000000 ;
			15'h000079BF : data <= 8'b00000000 ;
			15'h000079C0 : data <= 8'b00000000 ;
			15'h000079C1 : data <= 8'b00000000 ;
			15'h000079C2 : data <= 8'b00000000 ;
			15'h000079C3 : data <= 8'b00000000 ;
			15'h000079C4 : data <= 8'b00000000 ;
			15'h000079C5 : data <= 8'b00000000 ;
			15'h000079C6 : data <= 8'b00000000 ;
			15'h000079C7 : data <= 8'b00000000 ;
			15'h000079C8 : data <= 8'b00000000 ;
			15'h000079C9 : data <= 8'b00000000 ;
			15'h000079CA : data <= 8'b00000000 ;
			15'h000079CB : data <= 8'b00000000 ;
			15'h000079CC : data <= 8'b00000000 ;
			15'h000079CD : data <= 8'b00000000 ;
			15'h000079CE : data <= 8'b00000000 ;
			15'h000079CF : data <= 8'b00000000 ;
			15'h000079D0 : data <= 8'b00000000 ;
			15'h000079D1 : data <= 8'b00000000 ;
			15'h000079D2 : data <= 8'b00000000 ;
			15'h000079D3 : data <= 8'b00000000 ;
			15'h000079D4 : data <= 8'b00000000 ;
			15'h000079D5 : data <= 8'b00000000 ;
			15'h000079D6 : data <= 8'b00000000 ;
			15'h000079D7 : data <= 8'b00000000 ;
			15'h000079D8 : data <= 8'b00000000 ;
			15'h000079D9 : data <= 8'b00000000 ;
			15'h000079DA : data <= 8'b00000000 ;
			15'h000079DB : data <= 8'b00000000 ;
			15'h000079DC : data <= 8'b00000000 ;
			15'h000079DD : data <= 8'b00000000 ;
			15'h000079DE : data <= 8'b00000000 ;
			15'h000079DF : data <= 8'b00000000 ;
			15'h000079E0 : data <= 8'b00000000 ;
			15'h000079E1 : data <= 8'b00000000 ;
			15'h000079E2 : data <= 8'b00000000 ;
			15'h000079E3 : data <= 8'b00000000 ;
			15'h000079E4 : data <= 8'b00000000 ;
			15'h000079E5 : data <= 8'b00000000 ;
			15'h000079E6 : data <= 8'b00000000 ;
			15'h000079E7 : data <= 8'b00000000 ;
			15'h000079E8 : data <= 8'b00000000 ;
			15'h000079E9 : data <= 8'b00000000 ;
			15'h000079EA : data <= 8'b00000000 ;
			15'h000079EB : data <= 8'b00000000 ;
			15'h000079EC : data <= 8'b00000000 ;
			15'h000079ED : data <= 8'b00000000 ;
			15'h000079EE : data <= 8'b00000000 ;
			15'h000079EF : data <= 8'b00000000 ;
			15'h000079F0 : data <= 8'b00000000 ;
			15'h000079F1 : data <= 8'b00000000 ;
			15'h000079F2 : data <= 8'b00000000 ;
			15'h000079F3 : data <= 8'b00000000 ;
			15'h000079F4 : data <= 8'b00000000 ;
			15'h000079F5 : data <= 8'b00000000 ;
			15'h000079F6 : data <= 8'b00000000 ;
			15'h000079F7 : data <= 8'b00000000 ;
			15'h000079F8 : data <= 8'b00000000 ;
			15'h000079F9 : data <= 8'b00000000 ;
			15'h000079FA : data <= 8'b00000000 ;
			15'h000079FB : data <= 8'b00000000 ;
			15'h000079FC : data <= 8'b00000000 ;
			15'h000079FD : data <= 8'b00000000 ;
			15'h000079FE : data <= 8'b00000000 ;
			15'h000079FF : data <= 8'b00000000 ;
			15'h00007A00 : data <= 8'b00000000 ;
			15'h00007A01 : data <= 8'b00000000 ;
			15'h00007A02 : data <= 8'b00000000 ;
			15'h00007A03 : data <= 8'b00000000 ;
			15'h00007A04 : data <= 8'b00000000 ;
			15'h00007A05 : data <= 8'b00000000 ;
			15'h00007A06 : data <= 8'b00000000 ;
			15'h00007A07 : data <= 8'b00000000 ;
			15'h00007A08 : data <= 8'b00000000 ;
			15'h00007A09 : data <= 8'b00000000 ;
			15'h00007A0A : data <= 8'b00000000 ;
			15'h00007A0B : data <= 8'b00000000 ;
			15'h00007A0C : data <= 8'b00000000 ;
			15'h00007A0D : data <= 8'b00000000 ;
			15'h00007A0E : data <= 8'b00000000 ;
			15'h00007A0F : data <= 8'b00000000 ;
			15'h00007A10 : data <= 8'b00000000 ;
			15'h00007A11 : data <= 8'b00000000 ;
			15'h00007A12 : data <= 8'b00000000 ;
			15'h00007A13 : data <= 8'b00000000 ;
			15'h00007A14 : data <= 8'b00000000 ;
			15'h00007A15 : data <= 8'b00000000 ;
			15'h00007A16 : data <= 8'b00000000 ;
			15'h00007A17 : data <= 8'b00000000 ;
			15'h00007A18 : data <= 8'b00000000 ;
			15'h00007A19 : data <= 8'b00000000 ;
			15'h00007A1A : data <= 8'b00000000 ;
			15'h00007A1B : data <= 8'b00000000 ;
			15'h00007A1C : data <= 8'b00000000 ;
			15'h00007A1D : data <= 8'b00000000 ;
			15'h00007A1E : data <= 8'b00000000 ;
			15'h00007A1F : data <= 8'b00000000 ;
			15'h00007A20 : data <= 8'b00000000 ;
			15'h00007A21 : data <= 8'b00000000 ;
			15'h00007A22 : data <= 8'b00000000 ;
			15'h00007A23 : data <= 8'b00000000 ;
			15'h00007A24 : data <= 8'b00000000 ;
			15'h00007A25 : data <= 8'b00000000 ;
			15'h00007A26 : data <= 8'b00000000 ;
			15'h00007A27 : data <= 8'b00000000 ;
			15'h00007A28 : data <= 8'b00000000 ;
			15'h00007A29 : data <= 8'b00000000 ;
			15'h00007A2A : data <= 8'b00000000 ;
			15'h00007A2B : data <= 8'b00000000 ;
			15'h00007A2C : data <= 8'b00000000 ;
			15'h00007A2D : data <= 8'b00000000 ;
			15'h00007A2E : data <= 8'b00000000 ;
			15'h00007A2F : data <= 8'b00000000 ;
			15'h00007A30 : data <= 8'b00000000 ;
			15'h00007A31 : data <= 8'b00000000 ;
			15'h00007A32 : data <= 8'b00000000 ;
			15'h00007A33 : data <= 8'b00000000 ;
			15'h00007A34 : data <= 8'b00000000 ;
			15'h00007A35 : data <= 8'b00000000 ;
			15'h00007A36 : data <= 8'b00000000 ;
			15'h00007A37 : data <= 8'b00000000 ;
			15'h00007A38 : data <= 8'b00000000 ;
			15'h00007A39 : data <= 8'b00000000 ;
			15'h00007A3A : data <= 8'b00000000 ;
			15'h00007A3B : data <= 8'b00000000 ;
			15'h00007A3C : data <= 8'b00000000 ;
			15'h00007A3D : data <= 8'b00000000 ;
			15'h00007A3E : data <= 8'b00000000 ;
			15'h00007A3F : data <= 8'b00000000 ;
			15'h00007A40 : data <= 8'b00000000 ;
			15'h00007A41 : data <= 8'b00000000 ;
			15'h00007A42 : data <= 8'b00000000 ;
			15'h00007A43 : data <= 8'b00000000 ;
			15'h00007A44 : data <= 8'b00000000 ;
			15'h00007A45 : data <= 8'b00000000 ;
			15'h00007A46 : data <= 8'b00000000 ;
			15'h00007A47 : data <= 8'b00000000 ;
			15'h00007A48 : data <= 8'b00000000 ;
			15'h00007A49 : data <= 8'b00000000 ;
			15'h00007A4A : data <= 8'b00000000 ;
			15'h00007A4B : data <= 8'b00000000 ;
			15'h00007A4C : data <= 8'b00000000 ;
			15'h00007A4D : data <= 8'b00000000 ;
			15'h00007A4E : data <= 8'b00000000 ;
			15'h00007A4F : data <= 8'b00000000 ;
			15'h00007A50 : data <= 8'b00000000 ;
			15'h00007A51 : data <= 8'b00000000 ;
			15'h00007A52 : data <= 8'b00000000 ;
			15'h00007A53 : data <= 8'b00000000 ;
			15'h00007A54 : data <= 8'b00000000 ;
			15'h00007A55 : data <= 8'b00000000 ;
			15'h00007A56 : data <= 8'b00000000 ;
			15'h00007A57 : data <= 8'b00000000 ;
			15'h00007A58 : data <= 8'b00000000 ;
			15'h00007A59 : data <= 8'b00000000 ;
			15'h00007A5A : data <= 8'b00000000 ;
			15'h00007A5B : data <= 8'b00000000 ;
			15'h00007A5C : data <= 8'b00000000 ;
			15'h00007A5D : data <= 8'b00000000 ;
			15'h00007A5E : data <= 8'b00000000 ;
			15'h00007A5F : data <= 8'b00000000 ;
			15'h00007A60 : data <= 8'b00000000 ;
			15'h00007A61 : data <= 8'b00000000 ;
			15'h00007A62 : data <= 8'b00000000 ;
			15'h00007A63 : data <= 8'b00000000 ;
			15'h00007A64 : data <= 8'b00000000 ;
			15'h00007A65 : data <= 8'b00000000 ;
			15'h00007A66 : data <= 8'b00000000 ;
			15'h00007A67 : data <= 8'b00000000 ;
			15'h00007A68 : data <= 8'b00000000 ;
			15'h00007A69 : data <= 8'b00000000 ;
			15'h00007A6A : data <= 8'b00000000 ;
			15'h00007A6B : data <= 8'b00000000 ;
			15'h00007A6C : data <= 8'b00000000 ;
			15'h00007A6D : data <= 8'b00000000 ;
			15'h00007A6E : data <= 8'b00000000 ;
			15'h00007A6F : data <= 8'b00000000 ;
			15'h00007A70 : data <= 8'b00000000 ;
			15'h00007A71 : data <= 8'b00000000 ;
			15'h00007A72 : data <= 8'b00000000 ;
			15'h00007A73 : data <= 8'b00000000 ;
			15'h00007A74 : data <= 8'b00000000 ;
			15'h00007A75 : data <= 8'b00000000 ;
			15'h00007A76 : data <= 8'b00000000 ;
			15'h00007A77 : data <= 8'b00000000 ;
			15'h00007A78 : data <= 8'b00000000 ;
			15'h00007A79 : data <= 8'b00000000 ;
			15'h00007A7A : data <= 8'b00000000 ;
			15'h00007A7B : data <= 8'b00000000 ;
			15'h00007A7C : data <= 8'b00000000 ;
			15'h00007A7D : data <= 8'b00000000 ;
			15'h00007A7E : data <= 8'b00000000 ;
			15'h00007A7F : data <= 8'b00000000 ;
			15'h00007A80 : data <= 8'b00000000 ;
			15'h00007A81 : data <= 8'b00000000 ;
			15'h00007A82 : data <= 8'b00000000 ;
			15'h00007A83 : data <= 8'b00000000 ;
			15'h00007A84 : data <= 8'b00000000 ;
			15'h00007A85 : data <= 8'b00000000 ;
			15'h00007A86 : data <= 8'b00000000 ;
			15'h00007A87 : data <= 8'b00000000 ;
			15'h00007A88 : data <= 8'b00000000 ;
			15'h00007A89 : data <= 8'b00000000 ;
			15'h00007A8A : data <= 8'b00000000 ;
			15'h00007A8B : data <= 8'b00000000 ;
			15'h00007A8C : data <= 8'b00000000 ;
			15'h00007A8D : data <= 8'b00000000 ;
			15'h00007A8E : data <= 8'b00000000 ;
			15'h00007A8F : data <= 8'b00000000 ;
			15'h00007A90 : data <= 8'b00000000 ;
			15'h00007A91 : data <= 8'b00000000 ;
			15'h00007A92 : data <= 8'b00000000 ;
			15'h00007A93 : data <= 8'b00000000 ;
			15'h00007A94 : data <= 8'b00000000 ;
			15'h00007A95 : data <= 8'b00000000 ;
			15'h00007A96 : data <= 8'b00000000 ;
			15'h00007A97 : data <= 8'b00000000 ;
			15'h00007A98 : data <= 8'b00000000 ;
			15'h00007A99 : data <= 8'b00000000 ;
			15'h00007A9A : data <= 8'b00000000 ;
			15'h00007A9B : data <= 8'b00000000 ;
			15'h00007A9C : data <= 8'b00000000 ;
			15'h00007A9D : data <= 8'b00000000 ;
			15'h00007A9E : data <= 8'b00000000 ;
			15'h00007A9F : data <= 8'b00000000 ;
			15'h00007AA0 : data <= 8'b00000000 ;
			15'h00007AA1 : data <= 8'b00000000 ;
			15'h00007AA2 : data <= 8'b00000000 ;
			15'h00007AA3 : data <= 8'b00000000 ;
			15'h00007AA4 : data <= 8'b00000000 ;
			15'h00007AA5 : data <= 8'b00000000 ;
			15'h00007AA6 : data <= 8'b00000000 ;
			15'h00007AA7 : data <= 8'b00000000 ;
			15'h00007AA8 : data <= 8'b00000000 ;
			15'h00007AA9 : data <= 8'b00000000 ;
			15'h00007AAA : data <= 8'b00000000 ;
			15'h00007AAB : data <= 8'b00000000 ;
			15'h00007AAC : data <= 8'b00000000 ;
			15'h00007AAD : data <= 8'b00000000 ;
			15'h00007AAE : data <= 8'b00000000 ;
			15'h00007AAF : data <= 8'b00000000 ;
			15'h00007AB0 : data <= 8'b00000000 ;
			15'h00007AB1 : data <= 8'b00000000 ;
			15'h00007AB2 : data <= 8'b00000000 ;
			15'h00007AB3 : data <= 8'b00000000 ;
			15'h00007AB4 : data <= 8'b00000000 ;
			15'h00007AB5 : data <= 8'b00000000 ;
			15'h00007AB6 : data <= 8'b00000000 ;
			15'h00007AB7 : data <= 8'b00000000 ;
			15'h00007AB8 : data <= 8'b00000000 ;
			15'h00007AB9 : data <= 8'b00000000 ;
			15'h00007ABA : data <= 8'b00000000 ;
			15'h00007ABB : data <= 8'b00000000 ;
			15'h00007ABC : data <= 8'b00000000 ;
			15'h00007ABD : data <= 8'b00000000 ;
			15'h00007ABE : data <= 8'b00000000 ;
			15'h00007ABF : data <= 8'b00000000 ;
			15'h00007AC0 : data <= 8'b00000000 ;
			15'h00007AC1 : data <= 8'b00000000 ;
			15'h00007AC2 : data <= 8'b00000000 ;
			15'h00007AC3 : data <= 8'b00000000 ;
			15'h00007AC4 : data <= 8'b00000000 ;
			15'h00007AC5 : data <= 8'b00000000 ;
			15'h00007AC6 : data <= 8'b00000000 ;
			15'h00007AC7 : data <= 8'b00000000 ;
			15'h00007AC8 : data <= 8'b00000000 ;
			15'h00007AC9 : data <= 8'b00000000 ;
			15'h00007ACA : data <= 8'b00000000 ;
			15'h00007ACB : data <= 8'b00000000 ;
			15'h00007ACC : data <= 8'b00000000 ;
			15'h00007ACD : data <= 8'b00000000 ;
			15'h00007ACE : data <= 8'b00000000 ;
			15'h00007ACF : data <= 8'b00000000 ;
			15'h00007AD0 : data <= 8'b00000000 ;
			15'h00007AD1 : data <= 8'b00000000 ;
			15'h00007AD2 : data <= 8'b00000000 ;
			15'h00007AD3 : data <= 8'b00000000 ;
			15'h00007AD4 : data <= 8'b00000000 ;
			15'h00007AD5 : data <= 8'b00000000 ;
			15'h00007AD6 : data <= 8'b00000000 ;
			15'h00007AD7 : data <= 8'b00000000 ;
			15'h00007AD8 : data <= 8'b00000000 ;
			15'h00007AD9 : data <= 8'b00000000 ;
			15'h00007ADA : data <= 8'b00000000 ;
			15'h00007ADB : data <= 8'b00000000 ;
			15'h00007ADC : data <= 8'b00000000 ;
			15'h00007ADD : data <= 8'b00000000 ;
			15'h00007ADE : data <= 8'b00000000 ;
			15'h00007ADF : data <= 8'b00000000 ;
			15'h00007AE0 : data <= 8'b00000000 ;
			15'h00007AE1 : data <= 8'b00000000 ;
			15'h00007AE2 : data <= 8'b00000000 ;
			15'h00007AE3 : data <= 8'b00000000 ;
			15'h00007AE4 : data <= 8'b00000000 ;
			15'h00007AE5 : data <= 8'b00000000 ;
			15'h00007AE6 : data <= 8'b00000000 ;
			15'h00007AE7 : data <= 8'b00000000 ;
			15'h00007AE8 : data <= 8'b00000000 ;
			15'h00007AE9 : data <= 8'b00000000 ;
			15'h00007AEA : data <= 8'b00000000 ;
			15'h00007AEB : data <= 8'b00000000 ;
			15'h00007AEC : data <= 8'b00000000 ;
			15'h00007AED : data <= 8'b00000000 ;
			15'h00007AEE : data <= 8'b00000000 ;
			15'h00007AEF : data <= 8'b00000000 ;
			15'h00007AF0 : data <= 8'b00000000 ;
			15'h00007AF1 : data <= 8'b00000000 ;
			15'h00007AF2 : data <= 8'b00000000 ;
			15'h00007AF3 : data <= 8'b00000000 ;
			15'h00007AF4 : data <= 8'b00000000 ;
			15'h00007AF5 : data <= 8'b00000000 ;
			15'h00007AF6 : data <= 8'b00000000 ;
			15'h00007AF7 : data <= 8'b00000000 ;
			15'h00007AF8 : data <= 8'b00000000 ;
			15'h00007AF9 : data <= 8'b00000000 ;
			15'h00007AFA : data <= 8'b00000000 ;
			15'h00007AFB : data <= 8'b00000000 ;
			15'h00007AFC : data <= 8'b00000000 ;
			15'h00007AFD : data <= 8'b00000000 ;
			15'h00007AFE : data <= 8'b00000000 ;
			15'h00007AFF : data <= 8'b00000000 ;
			15'h00007B00 : data <= 8'b00000000 ;
			15'h00007B01 : data <= 8'b00000000 ;
			15'h00007B02 : data <= 8'b00000000 ;
			15'h00007B03 : data <= 8'b00000000 ;
			15'h00007B04 : data <= 8'b00000000 ;
			15'h00007B05 : data <= 8'b00000000 ;
			15'h00007B06 : data <= 8'b00000000 ;
			15'h00007B07 : data <= 8'b00000000 ;
			15'h00007B08 : data <= 8'b00000000 ;
			15'h00007B09 : data <= 8'b00000000 ;
			15'h00007B0A : data <= 8'b00000000 ;
			15'h00007B0B : data <= 8'b00000000 ;
			15'h00007B0C : data <= 8'b00000000 ;
			15'h00007B0D : data <= 8'b00000000 ;
			15'h00007B0E : data <= 8'b00000000 ;
			15'h00007B0F : data <= 8'b00000000 ;
			15'h00007B10 : data <= 8'b00000000 ;
			15'h00007B11 : data <= 8'b00000000 ;
			15'h00007B12 : data <= 8'b00000000 ;
			15'h00007B13 : data <= 8'b00000000 ;
			15'h00007B14 : data <= 8'b00000000 ;
			15'h00007B15 : data <= 8'b00000000 ;
			15'h00007B16 : data <= 8'b00000000 ;
			15'h00007B17 : data <= 8'b00000000 ;
			15'h00007B18 : data <= 8'b00000000 ;
			15'h00007B19 : data <= 8'b00000000 ;
			15'h00007B1A : data <= 8'b00000000 ;
			15'h00007B1B : data <= 8'b00000000 ;
			15'h00007B1C : data <= 8'b00000000 ;
			15'h00007B1D : data <= 8'b00000000 ;
			15'h00007B1E : data <= 8'b00000000 ;
			15'h00007B1F : data <= 8'b00000000 ;
			15'h00007B20 : data <= 8'b00000000 ;
			15'h00007B21 : data <= 8'b00000000 ;
			15'h00007B22 : data <= 8'b00000000 ;
			15'h00007B23 : data <= 8'b00000000 ;
			15'h00007B24 : data <= 8'b00000000 ;
			15'h00007B25 : data <= 8'b00000000 ;
			15'h00007B26 : data <= 8'b00000000 ;
			15'h00007B27 : data <= 8'b00000000 ;
			15'h00007B28 : data <= 8'b00000000 ;
			15'h00007B29 : data <= 8'b00000000 ;
			15'h00007B2A : data <= 8'b00000000 ;
			15'h00007B2B : data <= 8'b00000000 ;
			15'h00007B2C : data <= 8'b00000000 ;
			15'h00007B2D : data <= 8'b00000000 ;
			15'h00007B2E : data <= 8'b00000000 ;
			15'h00007B2F : data <= 8'b00000000 ;
			15'h00007B30 : data <= 8'b00000000 ;
			15'h00007B31 : data <= 8'b00000000 ;
			15'h00007B32 : data <= 8'b00000000 ;
			15'h00007B33 : data <= 8'b00000000 ;
			15'h00007B34 : data <= 8'b00000000 ;
			15'h00007B35 : data <= 8'b00000000 ;
			15'h00007B36 : data <= 8'b00000000 ;
			15'h00007B37 : data <= 8'b00000000 ;
			15'h00007B38 : data <= 8'b00000000 ;
			15'h00007B39 : data <= 8'b00000000 ;
			15'h00007B3A : data <= 8'b00000000 ;
			15'h00007B3B : data <= 8'b00000000 ;
			15'h00007B3C : data <= 8'b00000000 ;
			15'h00007B3D : data <= 8'b00000000 ;
			15'h00007B3E : data <= 8'b00000000 ;
			15'h00007B3F : data <= 8'b00000000 ;
			15'h00007B40 : data <= 8'b00000000 ;
			15'h00007B41 : data <= 8'b00000000 ;
			15'h00007B42 : data <= 8'b00000000 ;
			15'h00007B43 : data <= 8'b00000000 ;
			15'h00007B44 : data <= 8'b00000000 ;
			15'h00007B45 : data <= 8'b00000000 ;
			15'h00007B46 : data <= 8'b00000000 ;
			15'h00007B47 : data <= 8'b00000000 ;
			15'h00007B48 : data <= 8'b00000000 ;
			15'h00007B49 : data <= 8'b00000000 ;
			15'h00007B4A : data <= 8'b00000000 ;
			15'h00007B4B : data <= 8'b00000000 ;
			15'h00007B4C : data <= 8'b00000000 ;
			15'h00007B4D : data <= 8'b00000000 ;
			15'h00007B4E : data <= 8'b00000000 ;
			15'h00007B4F : data <= 8'b00000000 ;
			15'h00007B50 : data <= 8'b00000000 ;
			15'h00007B51 : data <= 8'b00000000 ;
			15'h00007B52 : data <= 8'b00000000 ;
			15'h00007B53 : data <= 8'b00000000 ;
			15'h00007B54 : data <= 8'b00000000 ;
			15'h00007B55 : data <= 8'b00000000 ;
			15'h00007B56 : data <= 8'b00000000 ;
			15'h00007B57 : data <= 8'b00000000 ;
			15'h00007B58 : data <= 8'b00000000 ;
			15'h00007B59 : data <= 8'b00000000 ;
			15'h00007B5A : data <= 8'b00000000 ;
			15'h00007B5B : data <= 8'b00000000 ;
			15'h00007B5C : data <= 8'b00000000 ;
			15'h00007B5D : data <= 8'b00000000 ;
			15'h00007B5E : data <= 8'b00000000 ;
			15'h00007B5F : data <= 8'b00000000 ;
			15'h00007B60 : data <= 8'b00000000 ;
			15'h00007B61 : data <= 8'b00000000 ;
			15'h00007B62 : data <= 8'b00000000 ;
			15'h00007B63 : data <= 8'b00000000 ;
			15'h00007B64 : data <= 8'b00000000 ;
			15'h00007B65 : data <= 8'b00000000 ;
			15'h00007B66 : data <= 8'b00000000 ;
			15'h00007B67 : data <= 8'b00000000 ;
			15'h00007B68 : data <= 8'b00000000 ;
			15'h00007B69 : data <= 8'b00000000 ;
			15'h00007B6A : data <= 8'b00000000 ;
			15'h00007B6B : data <= 8'b00000000 ;
			15'h00007B6C : data <= 8'b00000000 ;
			15'h00007B6D : data <= 8'b00000000 ;
			15'h00007B6E : data <= 8'b00000000 ;
			15'h00007B6F : data <= 8'b00000000 ;
			15'h00007B70 : data <= 8'b00000000 ;
			15'h00007B71 : data <= 8'b00000000 ;
			15'h00007B72 : data <= 8'b00000000 ;
			15'h00007B73 : data <= 8'b00000000 ;
			15'h00007B74 : data <= 8'b00000000 ;
			15'h00007B75 : data <= 8'b00000000 ;
			15'h00007B76 : data <= 8'b00000000 ;
			15'h00007B77 : data <= 8'b00000000 ;
			15'h00007B78 : data <= 8'b00000000 ;
			15'h00007B79 : data <= 8'b00000000 ;
			15'h00007B7A : data <= 8'b00000000 ;
			15'h00007B7B : data <= 8'b00000000 ;
			15'h00007B7C : data <= 8'b00000000 ;
			15'h00007B7D : data <= 8'b00000000 ;
			15'h00007B7E : data <= 8'b00000000 ;
			15'h00007B7F : data <= 8'b00000000 ;
			15'h00007B80 : data <= 8'b00000000 ;
			15'h00007B81 : data <= 8'b00000000 ;
			15'h00007B82 : data <= 8'b00000000 ;
			15'h00007B83 : data <= 8'b00000000 ;
			15'h00007B84 : data <= 8'b00000000 ;
			15'h00007B85 : data <= 8'b00000000 ;
			15'h00007B86 : data <= 8'b00000000 ;
			15'h00007B87 : data <= 8'b00000000 ;
			15'h00007B88 : data <= 8'b00000000 ;
			15'h00007B89 : data <= 8'b00000000 ;
			15'h00007B8A : data <= 8'b00000000 ;
			15'h00007B8B : data <= 8'b00000000 ;
			15'h00007B8C : data <= 8'b00000000 ;
			15'h00007B8D : data <= 8'b00000000 ;
			15'h00007B8E : data <= 8'b00000000 ;
			15'h00007B8F : data <= 8'b00000000 ;
			15'h00007B90 : data <= 8'b00000000 ;
			15'h00007B91 : data <= 8'b00000000 ;
			15'h00007B92 : data <= 8'b00000000 ;
			15'h00007B93 : data <= 8'b00000000 ;
			15'h00007B94 : data <= 8'b00000000 ;
			15'h00007B95 : data <= 8'b00000000 ;
			15'h00007B96 : data <= 8'b00000000 ;
			15'h00007B97 : data <= 8'b00000000 ;
			15'h00007B98 : data <= 8'b00000000 ;
			15'h00007B99 : data <= 8'b00000000 ;
			15'h00007B9A : data <= 8'b00000000 ;
			15'h00007B9B : data <= 8'b00000000 ;
			15'h00007B9C : data <= 8'b00000000 ;
			15'h00007B9D : data <= 8'b00000000 ;
			15'h00007B9E : data <= 8'b00000000 ;
			15'h00007B9F : data <= 8'b00000000 ;
			15'h00007BA0 : data <= 8'b00000000 ;
			15'h00007BA1 : data <= 8'b00000000 ;
			15'h00007BA2 : data <= 8'b00000000 ;
			15'h00007BA3 : data <= 8'b00000000 ;
			15'h00007BA4 : data <= 8'b00000000 ;
			15'h00007BA5 : data <= 8'b00000000 ;
			15'h00007BA6 : data <= 8'b00000000 ;
			15'h00007BA7 : data <= 8'b00000000 ;
			15'h00007BA8 : data <= 8'b00000000 ;
			15'h00007BA9 : data <= 8'b00000000 ;
			15'h00007BAA : data <= 8'b00000000 ;
			15'h00007BAB : data <= 8'b00000000 ;
			15'h00007BAC : data <= 8'b00000000 ;
			15'h00007BAD : data <= 8'b00000000 ;
			15'h00007BAE : data <= 8'b00000000 ;
			15'h00007BAF : data <= 8'b00000000 ;
			15'h00007BB0 : data <= 8'b00000000 ;
			15'h00007BB1 : data <= 8'b00000000 ;
			15'h00007BB2 : data <= 8'b00000000 ;
			15'h00007BB3 : data <= 8'b00000000 ;
			15'h00007BB4 : data <= 8'b00000000 ;
			15'h00007BB5 : data <= 8'b00000000 ;
			15'h00007BB6 : data <= 8'b00000000 ;
			15'h00007BB7 : data <= 8'b00000000 ;
			15'h00007BB8 : data <= 8'b00000000 ;
			15'h00007BB9 : data <= 8'b00000000 ;
			15'h00007BBA : data <= 8'b00000000 ;
			15'h00007BBB : data <= 8'b00000000 ;
			15'h00007BBC : data <= 8'b00000000 ;
			15'h00007BBD : data <= 8'b00000000 ;
			15'h00007BBE : data <= 8'b00000000 ;
			15'h00007BBF : data <= 8'b00000000 ;
			15'h00007BC0 : data <= 8'b00000000 ;
			15'h00007BC1 : data <= 8'b00000000 ;
			15'h00007BC2 : data <= 8'b00000000 ;
			15'h00007BC3 : data <= 8'b00000000 ;
			15'h00007BC4 : data <= 8'b00000000 ;
			15'h00007BC5 : data <= 8'b00000000 ;
			15'h00007BC6 : data <= 8'b00000000 ;
			15'h00007BC7 : data <= 8'b00000000 ;
			15'h00007BC8 : data <= 8'b00000000 ;
			15'h00007BC9 : data <= 8'b00000000 ;
			15'h00007BCA : data <= 8'b00000000 ;
			15'h00007BCB : data <= 8'b00000000 ;
			15'h00007BCC : data <= 8'b00000000 ;
			15'h00007BCD : data <= 8'b00000000 ;
			15'h00007BCE : data <= 8'b00000000 ;
			15'h00007BCF : data <= 8'b00000000 ;
			15'h00007BD0 : data <= 8'b00000000 ;
			15'h00007BD1 : data <= 8'b00000000 ;
			15'h00007BD2 : data <= 8'b00000000 ;
			15'h00007BD3 : data <= 8'b00000000 ;
			15'h00007BD4 : data <= 8'b00000000 ;
			15'h00007BD5 : data <= 8'b00000000 ;
			15'h00007BD6 : data <= 8'b00000000 ;
			15'h00007BD7 : data <= 8'b00000000 ;
			15'h00007BD8 : data <= 8'b00000000 ;
			15'h00007BD9 : data <= 8'b00000000 ;
			15'h00007BDA : data <= 8'b00000000 ;
			15'h00007BDB : data <= 8'b00000000 ;
			15'h00007BDC : data <= 8'b00000000 ;
			15'h00007BDD : data <= 8'b00000000 ;
			15'h00007BDE : data <= 8'b00000000 ;
			15'h00007BDF : data <= 8'b00000000 ;
			15'h00007BE0 : data <= 8'b00000000 ;
			15'h00007BE1 : data <= 8'b00000000 ;
			15'h00007BE2 : data <= 8'b00000000 ;
			15'h00007BE3 : data <= 8'b00000000 ;
			15'h00007BE4 : data <= 8'b00000000 ;
			15'h00007BE5 : data <= 8'b00000000 ;
			15'h00007BE6 : data <= 8'b00000000 ;
			15'h00007BE7 : data <= 8'b00000000 ;
			15'h00007BE8 : data <= 8'b00000000 ;
			15'h00007BE9 : data <= 8'b00000000 ;
			15'h00007BEA : data <= 8'b00000000 ;
			15'h00007BEB : data <= 8'b00000000 ;
			15'h00007BEC : data <= 8'b00000000 ;
			15'h00007BED : data <= 8'b00000000 ;
			15'h00007BEE : data <= 8'b00000000 ;
			15'h00007BEF : data <= 8'b00000000 ;
			15'h00007BF0 : data <= 8'b00000000 ;
			15'h00007BF1 : data <= 8'b00000000 ;
			15'h00007BF2 : data <= 8'b00000000 ;
			15'h00007BF3 : data <= 8'b00000000 ;
			15'h00007BF4 : data <= 8'b00000000 ;
			15'h00007BF5 : data <= 8'b00000000 ;
			15'h00007BF6 : data <= 8'b00000000 ;
			15'h00007BF7 : data <= 8'b00000000 ;
			15'h00007BF8 : data <= 8'b00000000 ;
			15'h00007BF9 : data <= 8'b00000000 ;
			15'h00007BFA : data <= 8'b00000000 ;
			15'h00007BFB : data <= 8'b00000000 ;
			15'h00007BFC : data <= 8'b00000000 ;
			15'h00007BFD : data <= 8'b00000000 ;
			15'h00007BFE : data <= 8'b00000000 ;
			15'h00007BFF : data <= 8'b00000000 ;
			15'h00007C00 : data <= 8'b00000000 ;
			15'h00007C01 : data <= 8'b00000000 ;
			15'h00007C02 : data <= 8'b00000000 ;
			15'h00007C03 : data <= 8'b00000000 ;
			15'h00007C04 : data <= 8'b00000000 ;
			15'h00007C05 : data <= 8'b00000000 ;
			15'h00007C06 : data <= 8'b00000000 ;
			15'h00007C07 : data <= 8'b00000000 ;
			15'h00007C08 : data <= 8'b00000000 ;
			15'h00007C09 : data <= 8'b00000000 ;
			15'h00007C0A : data <= 8'b00000000 ;
			15'h00007C0B : data <= 8'b00000000 ;
			15'h00007C0C : data <= 8'b00000000 ;
			15'h00007C0D : data <= 8'b00000000 ;
			15'h00007C0E : data <= 8'b00000000 ;
			15'h00007C0F : data <= 8'b00000000 ;
			15'h00007C10 : data <= 8'b00000000 ;
			15'h00007C11 : data <= 8'b00000000 ;
			15'h00007C12 : data <= 8'b00000000 ;
			15'h00007C13 : data <= 8'b00000000 ;
			15'h00007C14 : data <= 8'b00000000 ;
			15'h00007C15 : data <= 8'b00000000 ;
			15'h00007C16 : data <= 8'b00000000 ;
			15'h00007C17 : data <= 8'b00000000 ;
			15'h00007C18 : data <= 8'b00000000 ;
			15'h00007C19 : data <= 8'b00000000 ;
			15'h00007C1A : data <= 8'b00000000 ;
			15'h00007C1B : data <= 8'b00000000 ;
			15'h00007C1C : data <= 8'b00000000 ;
			15'h00007C1D : data <= 8'b00000000 ;
			15'h00007C1E : data <= 8'b00000000 ;
			15'h00007C1F : data <= 8'b00000000 ;
			15'h00007C20 : data <= 8'b00000000 ;
			15'h00007C21 : data <= 8'b00000000 ;
			15'h00007C22 : data <= 8'b00000000 ;
			15'h00007C23 : data <= 8'b00000000 ;
			15'h00007C24 : data <= 8'b00000000 ;
			15'h00007C25 : data <= 8'b00000000 ;
			15'h00007C26 : data <= 8'b00000000 ;
			15'h00007C27 : data <= 8'b00000000 ;
			15'h00007C28 : data <= 8'b00000000 ;
			15'h00007C29 : data <= 8'b00000000 ;
			15'h00007C2A : data <= 8'b00000000 ;
			15'h00007C2B : data <= 8'b00000000 ;
			15'h00007C2C : data <= 8'b00000000 ;
			15'h00007C2D : data <= 8'b00000000 ;
			15'h00007C2E : data <= 8'b00000000 ;
			15'h00007C2F : data <= 8'b00000000 ;
			15'h00007C30 : data <= 8'b00000000 ;
			15'h00007C31 : data <= 8'b00000000 ;
			15'h00007C32 : data <= 8'b00000000 ;
			15'h00007C33 : data <= 8'b00000000 ;
			15'h00007C34 : data <= 8'b00000000 ;
			15'h00007C35 : data <= 8'b00000000 ;
			15'h00007C36 : data <= 8'b00000000 ;
			15'h00007C37 : data <= 8'b00000000 ;
			15'h00007C38 : data <= 8'b00000000 ;
			15'h00007C39 : data <= 8'b00000000 ;
			15'h00007C3A : data <= 8'b00000000 ;
			15'h00007C3B : data <= 8'b00000000 ;
			15'h00007C3C : data <= 8'b00000000 ;
			15'h00007C3D : data <= 8'b00000000 ;
			15'h00007C3E : data <= 8'b00000000 ;
			15'h00007C3F : data <= 8'b00000000 ;
			15'h00007C40 : data <= 8'b00000000 ;
			15'h00007C41 : data <= 8'b00000000 ;
			15'h00007C42 : data <= 8'b00000000 ;
			15'h00007C43 : data <= 8'b00000000 ;
			15'h00007C44 : data <= 8'b00000000 ;
			15'h00007C45 : data <= 8'b00000000 ;
			15'h00007C46 : data <= 8'b00000000 ;
			15'h00007C47 : data <= 8'b00000000 ;
			15'h00007C48 : data <= 8'b00000000 ;
			15'h00007C49 : data <= 8'b00000000 ;
			15'h00007C4A : data <= 8'b00000000 ;
			15'h00007C4B : data <= 8'b00000000 ;
			15'h00007C4C : data <= 8'b00000000 ;
			15'h00007C4D : data <= 8'b00000000 ;
			15'h00007C4E : data <= 8'b00000000 ;
			15'h00007C4F : data <= 8'b00000000 ;
			15'h00007C50 : data <= 8'b00000000 ;
			15'h00007C51 : data <= 8'b00000000 ;
			15'h00007C52 : data <= 8'b00000000 ;
			15'h00007C53 : data <= 8'b00000000 ;
			15'h00007C54 : data <= 8'b00000000 ;
			15'h00007C55 : data <= 8'b00000000 ;
			15'h00007C56 : data <= 8'b00000000 ;
			15'h00007C57 : data <= 8'b00000000 ;
			15'h00007C58 : data <= 8'b00000000 ;
			15'h00007C59 : data <= 8'b00000000 ;
			15'h00007C5A : data <= 8'b00000000 ;
			15'h00007C5B : data <= 8'b00000000 ;
			15'h00007C5C : data <= 8'b00000000 ;
			15'h00007C5D : data <= 8'b00000000 ;
			15'h00007C5E : data <= 8'b00000000 ;
			15'h00007C5F : data <= 8'b00000000 ;
			15'h00007C60 : data <= 8'b00000000 ;
			15'h00007C61 : data <= 8'b00000000 ;
			15'h00007C62 : data <= 8'b00000000 ;
			15'h00007C63 : data <= 8'b00000000 ;
			15'h00007C64 : data <= 8'b00000000 ;
			15'h00007C65 : data <= 8'b00000000 ;
			15'h00007C66 : data <= 8'b00000000 ;
			15'h00007C67 : data <= 8'b00000000 ;
			15'h00007C68 : data <= 8'b00000000 ;
			15'h00007C69 : data <= 8'b00000000 ;
			15'h00007C6A : data <= 8'b00000000 ;
			15'h00007C6B : data <= 8'b00000000 ;
			15'h00007C6C : data <= 8'b00000000 ;
			15'h00007C6D : data <= 8'b00000000 ;
			15'h00007C6E : data <= 8'b00000000 ;
			15'h00007C6F : data <= 8'b00000000 ;
			15'h00007C70 : data <= 8'b00000000 ;
			15'h00007C71 : data <= 8'b00000000 ;
			15'h00007C72 : data <= 8'b00000000 ;
			15'h00007C73 : data <= 8'b00000000 ;
			15'h00007C74 : data <= 8'b00000000 ;
			15'h00007C75 : data <= 8'b00000000 ;
			15'h00007C76 : data <= 8'b00000000 ;
			15'h00007C77 : data <= 8'b00000000 ;
			15'h00007C78 : data <= 8'b00000000 ;
			15'h00007C79 : data <= 8'b00000000 ;
			15'h00007C7A : data <= 8'b00000000 ;
			15'h00007C7B : data <= 8'b00000000 ;
			15'h00007C7C : data <= 8'b00000000 ;
			15'h00007C7D : data <= 8'b00000000 ;
			15'h00007C7E : data <= 8'b00000000 ;
			15'h00007C7F : data <= 8'b00000000 ;
			15'h00007C80 : data <= 8'b00000000 ;
			15'h00007C81 : data <= 8'b00000000 ;
			15'h00007C82 : data <= 8'b00000000 ;
			15'h00007C83 : data <= 8'b00000000 ;
			15'h00007C84 : data <= 8'b00000000 ;
			15'h00007C85 : data <= 8'b00000000 ;
			15'h00007C86 : data <= 8'b00000000 ;
			15'h00007C87 : data <= 8'b00000000 ;
			15'h00007C88 : data <= 8'b00000000 ;
			15'h00007C89 : data <= 8'b00000000 ;
			15'h00007C8A : data <= 8'b00000000 ;
			15'h00007C8B : data <= 8'b00000000 ;
			15'h00007C8C : data <= 8'b00000000 ;
			15'h00007C8D : data <= 8'b00000000 ;
			15'h00007C8E : data <= 8'b00000000 ;
			15'h00007C8F : data <= 8'b00000000 ;
			15'h00007C90 : data <= 8'b00000000 ;
			15'h00007C91 : data <= 8'b00000000 ;
			15'h00007C92 : data <= 8'b00000000 ;
			15'h00007C93 : data <= 8'b00000000 ;
			15'h00007C94 : data <= 8'b00000000 ;
			15'h00007C95 : data <= 8'b00000000 ;
			15'h00007C96 : data <= 8'b00000000 ;
			15'h00007C97 : data <= 8'b00000000 ;
			15'h00007C98 : data <= 8'b00000000 ;
			15'h00007C99 : data <= 8'b00000000 ;
			15'h00007C9A : data <= 8'b00000000 ;
			15'h00007C9B : data <= 8'b00000000 ;
			15'h00007C9C : data <= 8'b00000000 ;
			15'h00007C9D : data <= 8'b00000000 ;
			15'h00007C9E : data <= 8'b00000000 ;
			15'h00007C9F : data <= 8'b00000000 ;
			15'h00007CA0 : data <= 8'b00000000 ;
			15'h00007CA1 : data <= 8'b00000000 ;
			15'h00007CA2 : data <= 8'b00000000 ;
			15'h00007CA3 : data <= 8'b00000000 ;
			15'h00007CA4 : data <= 8'b00000000 ;
			15'h00007CA5 : data <= 8'b00000000 ;
			15'h00007CA6 : data <= 8'b00000000 ;
			15'h00007CA7 : data <= 8'b00000000 ;
			15'h00007CA8 : data <= 8'b00000000 ;
			15'h00007CA9 : data <= 8'b00000000 ;
			15'h00007CAA : data <= 8'b00000000 ;
			15'h00007CAB : data <= 8'b00000000 ;
			15'h00007CAC : data <= 8'b00000000 ;
			15'h00007CAD : data <= 8'b00000000 ;
			15'h00007CAE : data <= 8'b00000000 ;
			15'h00007CAF : data <= 8'b00000000 ;
			15'h00007CB0 : data <= 8'b00000000 ;
			15'h00007CB1 : data <= 8'b00000000 ;
			15'h00007CB2 : data <= 8'b00000000 ;
			15'h00007CB3 : data <= 8'b00000000 ;
			15'h00007CB4 : data <= 8'b00000000 ;
			15'h00007CB5 : data <= 8'b00000000 ;
			15'h00007CB6 : data <= 8'b00000000 ;
			15'h00007CB7 : data <= 8'b00000000 ;
			15'h00007CB8 : data <= 8'b00000000 ;
			15'h00007CB9 : data <= 8'b00000000 ;
			15'h00007CBA : data <= 8'b00000000 ;
			15'h00007CBB : data <= 8'b00000000 ;
			15'h00007CBC : data <= 8'b00000000 ;
			15'h00007CBD : data <= 8'b00000000 ;
			15'h00007CBE : data <= 8'b00000000 ;
			15'h00007CBF : data <= 8'b00000000 ;
			15'h00007CC0 : data <= 8'b00000000 ;
			15'h00007CC1 : data <= 8'b00000000 ;
			15'h00007CC2 : data <= 8'b00000000 ;
			15'h00007CC3 : data <= 8'b00000000 ;
			15'h00007CC4 : data <= 8'b00000000 ;
			15'h00007CC5 : data <= 8'b00000000 ;
			15'h00007CC6 : data <= 8'b00000000 ;
			15'h00007CC7 : data <= 8'b00000000 ;
			15'h00007CC8 : data <= 8'b00000000 ;
			15'h00007CC9 : data <= 8'b00000000 ;
			15'h00007CCA : data <= 8'b00000000 ;
			15'h00007CCB : data <= 8'b00000000 ;
			15'h00007CCC : data <= 8'b00000000 ;
			15'h00007CCD : data <= 8'b00000000 ;
			15'h00007CCE : data <= 8'b00000000 ;
			15'h00007CCF : data <= 8'b00000000 ;
			15'h00007CD0 : data <= 8'b00000000 ;
			15'h00007CD1 : data <= 8'b00000000 ;
			15'h00007CD2 : data <= 8'b00000000 ;
			15'h00007CD3 : data <= 8'b00000000 ;
			15'h00007CD4 : data <= 8'b00000000 ;
			15'h00007CD5 : data <= 8'b00000000 ;
			15'h00007CD6 : data <= 8'b00000000 ;
			15'h00007CD7 : data <= 8'b00000000 ;
			15'h00007CD8 : data <= 8'b00000000 ;
			15'h00007CD9 : data <= 8'b00000000 ;
			15'h00007CDA : data <= 8'b00000000 ;
			15'h00007CDB : data <= 8'b00000000 ;
			15'h00007CDC : data <= 8'b00000000 ;
			15'h00007CDD : data <= 8'b00000000 ;
			15'h00007CDE : data <= 8'b00000000 ;
			15'h00007CDF : data <= 8'b00000000 ;
			15'h00007CE0 : data <= 8'b00000000 ;
			15'h00007CE1 : data <= 8'b00000000 ;
			15'h00007CE2 : data <= 8'b00000000 ;
			15'h00007CE3 : data <= 8'b00000000 ;
			15'h00007CE4 : data <= 8'b00000000 ;
			15'h00007CE5 : data <= 8'b00000000 ;
			15'h00007CE6 : data <= 8'b00000000 ;
			15'h00007CE7 : data <= 8'b00000000 ;
			15'h00007CE8 : data <= 8'b00000000 ;
			15'h00007CE9 : data <= 8'b00000000 ;
			15'h00007CEA : data <= 8'b00000000 ;
			15'h00007CEB : data <= 8'b00000000 ;
			15'h00007CEC : data <= 8'b00000000 ;
			15'h00007CED : data <= 8'b00000000 ;
			15'h00007CEE : data <= 8'b00000000 ;
			15'h00007CEF : data <= 8'b00000000 ;
			15'h00007CF0 : data <= 8'b00000000 ;
			15'h00007CF1 : data <= 8'b00000000 ;
			15'h00007CF2 : data <= 8'b00000000 ;
			15'h00007CF3 : data <= 8'b00000000 ;
			15'h00007CF4 : data <= 8'b00000000 ;
			15'h00007CF5 : data <= 8'b00000000 ;
			15'h00007CF6 : data <= 8'b00000000 ;
			15'h00007CF7 : data <= 8'b00000000 ;
			15'h00007CF8 : data <= 8'b00000000 ;
			15'h00007CF9 : data <= 8'b00000000 ;
			15'h00007CFA : data <= 8'b00000000 ;
			15'h00007CFB : data <= 8'b00000000 ;
			15'h00007CFC : data <= 8'b00000000 ;
			15'h00007CFD : data <= 8'b00000000 ;
			15'h00007CFE : data <= 8'b00000000 ;
			15'h00007CFF : data <= 8'b00000000 ;
			15'h00007D00 : data <= 8'b00000000 ;
			15'h00007D01 : data <= 8'b00000000 ;
			15'h00007D02 : data <= 8'b00000000 ;
			15'h00007D03 : data <= 8'b00000000 ;
			15'h00007D04 : data <= 8'b00000000 ;
			15'h00007D05 : data <= 8'b00000000 ;
			15'h00007D06 : data <= 8'b00000000 ;
			15'h00007D07 : data <= 8'b00000000 ;
			15'h00007D08 : data <= 8'b00000000 ;
			15'h00007D09 : data <= 8'b00000000 ;
			15'h00007D0A : data <= 8'b00000000 ;
			15'h00007D0B : data <= 8'b00000000 ;
			15'h00007D0C : data <= 8'b00000000 ;
			15'h00007D0D : data <= 8'b00000000 ;
			15'h00007D0E : data <= 8'b00000000 ;
			15'h00007D0F : data <= 8'b00000000 ;
			15'h00007D10 : data <= 8'b00000000 ;
			15'h00007D11 : data <= 8'b00000000 ;
			15'h00007D12 : data <= 8'b00000000 ;
			15'h00007D13 : data <= 8'b00000000 ;
			15'h00007D14 : data <= 8'b00000000 ;
			15'h00007D15 : data <= 8'b00000000 ;
			15'h00007D16 : data <= 8'b00000000 ;
			15'h00007D17 : data <= 8'b00000000 ;
			15'h00007D18 : data <= 8'b00000000 ;
			15'h00007D19 : data <= 8'b00000000 ;
			15'h00007D1A : data <= 8'b00000000 ;
			15'h00007D1B : data <= 8'b00000000 ;
			15'h00007D1C : data <= 8'b00000000 ;
			15'h00007D1D : data <= 8'b00000000 ;
			15'h00007D1E : data <= 8'b00000000 ;
			15'h00007D1F : data <= 8'b00000000 ;
			15'h00007D20 : data <= 8'b00000000 ;
			15'h00007D21 : data <= 8'b00000000 ;
			15'h00007D22 : data <= 8'b00000000 ;
			15'h00007D23 : data <= 8'b00000000 ;
			15'h00007D24 : data <= 8'b00000000 ;
			15'h00007D25 : data <= 8'b00000000 ;
			15'h00007D26 : data <= 8'b00000000 ;
			15'h00007D27 : data <= 8'b00000000 ;
			15'h00007D28 : data <= 8'b00000000 ;
			15'h00007D29 : data <= 8'b00000000 ;
			15'h00007D2A : data <= 8'b00000000 ;
			15'h00007D2B : data <= 8'b00000000 ;
			15'h00007D2C : data <= 8'b00000000 ;
			15'h00007D2D : data <= 8'b00000000 ;
			15'h00007D2E : data <= 8'b00000000 ;
			15'h00007D2F : data <= 8'b00000000 ;
			15'h00007D30 : data <= 8'b00000000 ;
			15'h00007D31 : data <= 8'b00000000 ;
			15'h00007D32 : data <= 8'b00000000 ;
			15'h00007D33 : data <= 8'b00000000 ;
			15'h00007D34 : data <= 8'b00000000 ;
			15'h00007D35 : data <= 8'b00000000 ;
			15'h00007D36 : data <= 8'b00000000 ;
			15'h00007D37 : data <= 8'b00000000 ;
			15'h00007D38 : data <= 8'b00000000 ;
			15'h00007D39 : data <= 8'b00000000 ;
			15'h00007D3A : data <= 8'b00000000 ;
			15'h00007D3B : data <= 8'b00000000 ;
			15'h00007D3C : data <= 8'b00000000 ;
			15'h00007D3D : data <= 8'b00000000 ;
			15'h00007D3E : data <= 8'b00000000 ;
			15'h00007D3F : data <= 8'b00000000 ;
			15'h00007D40 : data <= 8'b00000000 ;
			15'h00007D41 : data <= 8'b00000000 ;
			15'h00007D42 : data <= 8'b00000000 ;
			15'h00007D43 : data <= 8'b00000000 ;
			15'h00007D44 : data <= 8'b00000000 ;
			15'h00007D45 : data <= 8'b00000000 ;
			15'h00007D46 : data <= 8'b00000000 ;
			15'h00007D47 : data <= 8'b00000000 ;
			15'h00007D48 : data <= 8'b00000000 ;
			15'h00007D49 : data <= 8'b00000000 ;
			15'h00007D4A : data <= 8'b00000000 ;
			15'h00007D4B : data <= 8'b00000000 ;
			15'h00007D4C : data <= 8'b00000000 ;
			15'h00007D4D : data <= 8'b00000000 ;
			15'h00007D4E : data <= 8'b00000000 ;
			15'h00007D4F : data <= 8'b00000000 ;
			15'h00007D50 : data <= 8'b00000000 ;
			15'h00007D51 : data <= 8'b00000000 ;
			15'h00007D52 : data <= 8'b00000000 ;
			15'h00007D53 : data <= 8'b00000000 ;
			15'h00007D54 : data <= 8'b00000000 ;
			15'h00007D55 : data <= 8'b00000000 ;
			15'h00007D56 : data <= 8'b00000000 ;
			15'h00007D57 : data <= 8'b00000000 ;
			15'h00007D58 : data <= 8'b00000000 ;
			15'h00007D59 : data <= 8'b00000000 ;
			15'h00007D5A : data <= 8'b00000000 ;
			15'h00007D5B : data <= 8'b00000000 ;
			15'h00007D5C : data <= 8'b00000000 ;
			15'h00007D5D : data <= 8'b00000000 ;
			15'h00007D5E : data <= 8'b00000000 ;
			15'h00007D5F : data <= 8'b00000000 ;
			15'h00007D60 : data <= 8'b00000000 ;
			15'h00007D61 : data <= 8'b00000000 ;
			15'h00007D62 : data <= 8'b00000000 ;
			15'h00007D63 : data <= 8'b00000000 ;
			15'h00007D64 : data <= 8'b00000000 ;
			15'h00007D65 : data <= 8'b00000000 ;
			15'h00007D66 : data <= 8'b00000000 ;
			15'h00007D67 : data <= 8'b00000000 ;
			15'h00007D68 : data <= 8'b00000000 ;
			15'h00007D69 : data <= 8'b00000000 ;
			15'h00007D6A : data <= 8'b00000000 ;
			15'h00007D6B : data <= 8'b00000000 ;
			15'h00007D6C : data <= 8'b00000000 ;
			15'h00007D6D : data <= 8'b00000000 ;
			15'h00007D6E : data <= 8'b00000000 ;
			15'h00007D6F : data <= 8'b00000000 ;
			15'h00007D70 : data <= 8'b00000000 ;
			15'h00007D71 : data <= 8'b00000000 ;
			15'h00007D72 : data <= 8'b00000000 ;
			15'h00007D73 : data <= 8'b00000000 ;
			15'h00007D74 : data <= 8'b00000000 ;
			15'h00007D75 : data <= 8'b00000000 ;
			15'h00007D76 : data <= 8'b00000000 ;
			15'h00007D77 : data <= 8'b00000000 ;
			15'h00007D78 : data <= 8'b00000000 ;
			15'h00007D79 : data <= 8'b00000000 ;
			15'h00007D7A : data <= 8'b00000000 ;
			15'h00007D7B : data <= 8'b00000000 ;
			15'h00007D7C : data <= 8'b00000000 ;
			15'h00007D7D : data <= 8'b00000000 ;
			15'h00007D7E : data <= 8'b00000000 ;
			15'h00007D7F : data <= 8'b00000000 ;
			15'h00007D80 : data <= 8'b00000000 ;
			15'h00007D81 : data <= 8'b00000000 ;
			15'h00007D82 : data <= 8'b00000000 ;
			15'h00007D83 : data <= 8'b00000000 ;
			15'h00007D84 : data <= 8'b00000000 ;
			15'h00007D85 : data <= 8'b00000000 ;
			15'h00007D86 : data <= 8'b00000000 ;
			15'h00007D87 : data <= 8'b00000000 ;
			15'h00007D88 : data <= 8'b00000000 ;
			15'h00007D89 : data <= 8'b00000000 ;
			15'h00007D8A : data <= 8'b00000000 ;
			15'h00007D8B : data <= 8'b00000000 ;
			15'h00007D8C : data <= 8'b00000000 ;
			15'h00007D8D : data <= 8'b00000000 ;
			15'h00007D8E : data <= 8'b00000000 ;
			15'h00007D8F : data <= 8'b00000000 ;
			15'h00007D90 : data <= 8'b00000000 ;
			15'h00007D91 : data <= 8'b00000000 ;
			15'h00007D92 : data <= 8'b00000000 ;
			15'h00007D93 : data <= 8'b00000000 ;
			15'h00007D94 : data <= 8'b00000000 ;
			15'h00007D95 : data <= 8'b00000000 ;
			15'h00007D96 : data <= 8'b00000000 ;
			15'h00007D97 : data <= 8'b00000000 ;
			15'h00007D98 : data <= 8'b00000000 ;
			15'h00007D99 : data <= 8'b00000000 ;
			15'h00007D9A : data <= 8'b00000000 ;
			15'h00007D9B : data <= 8'b00000000 ;
			15'h00007D9C : data <= 8'b00000000 ;
			15'h00007D9D : data <= 8'b00000000 ;
			15'h00007D9E : data <= 8'b00000000 ;
			15'h00007D9F : data <= 8'b00000000 ;
			15'h00007DA0 : data <= 8'b00000000 ;
			15'h00007DA1 : data <= 8'b00000000 ;
			15'h00007DA2 : data <= 8'b00000000 ;
			15'h00007DA3 : data <= 8'b00000000 ;
			15'h00007DA4 : data <= 8'b00000000 ;
			15'h00007DA5 : data <= 8'b00000000 ;
			15'h00007DA6 : data <= 8'b00000000 ;
			15'h00007DA7 : data <= 8'b00000000 ;
			15'h00007DA8 : data <= 8'b00000000 ;
			15'h00007DA9 : data <= 8'b00000000 ;
			15'h00007DAA : data <= 8'b00000000 ;
			15'h00007DAB : data <= 8'b00000000 ;
			15'h00007DAC : data <= 8'b00000000 ;
			15'h00007DAD : data <= 8'b00000000 ;
			15'h00007DAE : data <= 8'b00000000 ;
			15'h00007DAF : data <= 8'b00000000 ;
			15'h00007DB0 : data <= 8'b00000000 ;
			15'h00007DB1 : data <= 8'b00000000 ;
			15'h00007DB2 : data <= 8'b00000000 ;
			15'h00007DB3 : data <= 8'b00000000 ;
			15'h00007DB4 : data <= 8'b00000000 ;
			15'h00007DB5 : data <= 8'b00000000 ;
			15'h00007DB6 : data <= 8'b00000000 ;
			15'h00007DB7 : data <= 8'b00000000 ;
			15'h00007DB8 : data <= 8'b00000000 ;
			15'h00007DB9 : data <= 8'b00000000 ;
			15'h00007DBA : data <= 8'b00000000 ;
			15'h00007DBB : data <= 8'b00000000 ;
			15'h00007DBC : data <= 8'b00000000 ;
			15'h00007DBD : data <= 8'b00000000 ;
			15'h00007DBE : data <= 8'b00000000 ;
			15'h00007DBF : data <= 8'b00000000 ;
			15'h00007DC0 : data <= 8'b00000000 ;
			15'h00007DC1 : data <= 8'b00000000 ;
			15'h00007DC2 : data <= 8'b00000000 ;
			15'h00007DC3 : data <= 8'b00000000 ;
			15'h00007DC4 : data <= 8'b00000000 ;
			15'h00007DC5 : data <= 8'b00000000 ;
			15'h00007DC6 : data <= 8'b00000000 ;
			15'h00007DC7 : data <= 8'b00000000 ;
			15'h00007DC8 : data <= 8'b00000000 ;
			15'h00007DC9 : data <= 8'b00000000 ;
			15'h00007DCA : data <= 8'b00000000 ;
			15'h00007DCB : data <= 8'b00000000 ;
			15'h00007DCC : data <= 8'b00000000 ;
			15'h00007DCD : data <= 8'b00000000 ;
			15'h00007DCE : data <= 8'b00000000 ;
			15'h00007DCF : data <= 8'b00000000 ;
			15'h00007DD0 : data <= 8'b00000000 ;
			15'h00007DD1 : data <= 8'b00000000 ;
			15'h00007DD2 : data <= 8'b00000000 ;
			15'h00007DD3 : data <= 8'b00000000 ;
			15'h00007DD4 : data <= 8'b00000000 ;
			15'h00007DD5 : data <= 8'b00000000 ;
			15'h00007DD6 : data <= 8'b00000000 ;
			15'h00007DD7 : data <= 8'b00000000 ;
			15'h00007DD8 : data <= 8'b00000000 ;
			15'h00007DD9 : data <= 8'b00000000 ;
			15'h00007DDA : data <= 8'b00000000 ;
			15'h00007DDB : data <= 8'b00000000 ;
			15'h00007DDC : data <= 8'b00000000 ;
			15'h00007DDD : data <= 8'b00000000 ;
			15'h00007DDE : data <= 8'b00000000 ;
			15'h00007DDF : data <= 8'b00000000 ;
			15'h00007DE0 : data <= 8'b00000000 ;
			15'h00007DE1 : data <= 8'b00000000 ;
			15'h00007DE2 : data <= 8'b00000000 ;
			15'h00007DE3 : data <= 8'b00000000 ;
			15'h00007DE4 : data <= 8'b00000000 ;
			15'h00007DE5 : data <= 8'b00000000 ;
			15'h00007DE6 : data <= 8'b00000000 ;
			15'h00007DE7 : data <= 8'b00000000 ;
			15'h00007DE8 : data <= 8'b00000000 ;
			15'h00007DE9 : data <= 8'b00000000 ;
			15'h00007DEA : data <= 8'b00000000 ;
			15'h00007DEB : data <= 8'b00000000 ;
			15'h00007DEC : data <= 8'b00000000 ;
			15'h00007DED : data <= 8'b00000000 ;
			15'h00007DEE : data <= 8'b00000000 ;
			15'h00007DEF : data <= 8'b00000000 ;
			15'h00007DF0 : data <= 8'b00000000 ;
			15'h00007DF1 : data <= 8'b00000000 ;
			15'h00007DF2 : data <= 8'b00000000 ;
			15'h00007DF3 : data <= 8'b00000000 ;
			15'h00007DF4 : data <= 8'b00000000 ;
			15'h00007DF5 : data <= 8'b00000000 ;
			15'h00007DF6 : data <= 8'b00000000 ;
			15'h00007DF7 : data <= 8'b00000000 ;
			15'h00007DF8 : data <= 8'b00000000 ;
			15'h00007DF9 : data <= 8'b00000000 ;
			15'h00007DFA : data <= 8'b00000000 ;
			15'h00007DFB : data <= 8'b00000000 ;
			15'h00007DFC : data <= 8'b00000000 ;
			15'h00007DFD : data <= 8'b00000000 ;
			15'h00007DFE : data <= 8'b00000000 ;
			15'h00007DFF : data <= 8'b00000000 ;
			15'h00007E00 : data <= 8'b00000000 ;
			15'h00007E01 : data <= 8'b00000000 ;
			15'h00007E02 : data <= 8'b00000000 ;
			15'h00007E03 : data <= 8'b00000000 ;
			15'h00007E04 : data <= 8'b00000000 ;
			15'h00007E05 : data <= 8'b00000000 ;
			15'h00007E06 : data <= 8'b00000000 ;
			15'h00007E07 : data <= 8'b00000000 ;
			15'h00007E08 : data <= 8'b00000000 ;
			15'h00007E09 : data <= 8'b00000000 ;
			15'h00007E0A : data <= 8'b00000000 ;
			15'h00007E0B : data <= 8'b00000000 ;
			15'h00007E0C : data <= 8'b00000000 ;
			15'h00007E0D : data <= 8'b00000000 ;
			15'h00007E0E : data <= 8'b00000000 ;
			15'h00007E0F : data <= 8'b00000000 ;
			15'h00007E10 : data <= 8'b00000000 ;
			15'h00007E11 : data <= 8'b00000000 ;
			15'h00007E12 : data <= 8'b00000000 ;
			15'h00007E13 : data <= 8'b00000000 ;
			15'h00007E14 : data <= 8'b00000000 ;
			15'h00007E15 : data <= 8'b00000000 ;
			15'h00007E16 : data <= 8'b00000000 ;
			15'h00007E17 : data <= 8'b00000000 ;
			15'h00007E18 : data <= 8'b00000000 ;
			15'h00007E19 : data <= 8'b00000000 ;
			15'h00007E1A : data <= 8'b00000000 ;
			15'h00007E1B : data <= 8'b00000000 ;
			15'h00007E1C : data <= 8'b00000000 ;
			15'h00007E1D : data <= 8'b00000000 ;
			15'h00007E1E : data <= 8'b00000000 ;
			15'h00007E1F : data <= 8'b00000000 ;
			15'h00007E20 : data <= 8'b00000000 ;
			15'h00007E21 : data <= 8'b00000000 ;
			15'h00007E22 : data <= 8'b00000000 ;
			15'h00007E23 : data <= 8'b00000000 ;
			15'h00007E24 : data <= 8'b00000000 ;
			15'h00007E25 : data <= 8'b00000000 ;
			15'h00007E26 : data <= 8'b00000000 ;
			15'h00007E27 : data <= 8'b00000000 ;
			15'h00007E28 : data <= 8'b00000000 ;
			15'h00007E29 : data <= 8'b00000000 ;
			15'h00007E2A : data <= 8'b00000000 ;
			15'h00007E2B : data <= 8'b00000000 ;
			15'h00007E2C : data <= 8'b00000000 ;
			15'h00007E2D : data <= 8'b00000000 ;
			15'h00007E2E : data <= 8'b00000000 ;
			15'h00007E2F : data <= 8'b00000000 ;
			15'h00007E30 : data <= 8'b00000000 ;
			15'h00007E31 : data <= 8'b00000000 ;
			15'h00007E32 : data <= 8'b00000000 ;
			15'h00007E33 : data <= 8'b00000000 ;
			15'h00007E34 : data <= 8'b00000000 ;
			15'h00007E35 : data <= 8'b00000000 ;
			15'h00007E36 : data <= 8'b00000000 ;
			15'h00007E37 : data <= 8'b00000000 ;
			15'h00007E38 : data <= 8'b00000000 ;
			15'h00007E39 : data <= 8'b00000000 ;
			15'h00007E3A : data <= 8'b00000000 ;
			15'h00007E3B : data <= 8'b00000000 ;
			15'h00007E3C : data <= 8'b00000000 ;
			15'h00007E3D : data <= 8'b00000000 ;
			15'h00007E3E : data <= 8'b00000000 ;
			15'h00007E3F : data <= 8'b00000000 ;
			15'h00007E40 : data <= 8'b00000000 ;
			15'h00007E41 : data <= 8'b00000000 ;
			15'h00007E42 : data <= 8'b00000000 ;
			15'h00007E43 : data <= 8'b00000000 ;
			15'h00007E44 : data <= 8'b00000000 ;
			15'h00007E45 : data <= 8'b00000000 ;
			15'h00007E46 : data <= 8'b00000000 ;
			15'h00007E47 : data <= 8'b00000000 ;
			15'h00007E48 : data <= 8'b00000000 ;
			15'h00007E49 : data <= 8'b00000000 ;
			15'h00007E4A : data <= 8'b00000000 ;
			15'h00007E4B : data <= 8'b00000000 ;
			15'h00007E4C : data <= 8'b00000000 ;
			15'h00007E4D : data <= 8'b00000000 ;
			15'h00007E4E : data <= 8'b00000000 ;
			15'h00007E4F : data <= 8'b00000000 ;
			15'h00007E50 : data <= 8'b00000000 ;
			15'h00007E51 : data <= 8'b00000000 ;
			15'h00007E52 : data <= 8'b00000000 ;
			15'h00007E53 : data <= 8'b00000000 ;
			15'h00007E54 : data <= 8'b00000000 ;
			15'h00007E55 : data <= 8'b00000000 ;
			15'h00007E56 : data <= 8'b00000000 ;
			15'h00007E57 : data <= 8'b00000000 ;
			15'h00007E58 : data <= 8'b00000000 ;
			15'h00007E59 : data <= 8'b00000000 ;
			15'h00007E5A : data <= 8'b00000000 ;
			15'h00007E5B : data <= 8'b00000000 ;
			15'h00007E5C : data <= 8'b00000000 ;
			15'h00007E5D : data <= 8'b00000000 ;
			15'h00007E5E : data <= 8'b00000000 ;
			15'h00007E5F : data <= 8'b00000000 ;
			15'h00007E60 : data <= 8'b00000000 ;
			15'h00007E61 : data <= 8'b00000000 ;
			15'h00007E62 : data <= 8'b00000000 ;
			15'h00007E63 : data <= 8'b00000000 ;
			15'h00007E64 : data <= 8'b00000000 ;
			15'h00007E65 : data <= 8'b00000000 ;
			15'h00007E66 : data <= 8'b00000000 ;
			15'h00007E67 : data <= 8'b00000000 ;
			15'h00007E68 : data <= 8'b00000000 ;
			15'h00007E69 : data <= 8'b00000000 ;
			15'h00007E6A : data <= 8'b00000000 ;
			15'h00007E6B : data <= 8'b00000000 ;
			15'h00007E6C : data <= 8'b00000000 ;
			15'h00007E6D : data <= 8'b00000000 ;
			15'h00007E6E : data <= 8'b00000000 ;
			15'h00007E6F : data <= 8'b00000000 ;
			15'h00007E70 : data <= 8'b00000000 ;
			15'h00007E71 : data <= 8'b00000000 ;
			15'h00007E72 : data <= 8'b00000000 ;
			15'h00007E73 : data <= 8'b00000000 ;
			15'h00007E74 : data <= 8'b00000000 ;
			15'h00007E75 : data <= 8'b00000000 ;
			15'h00007E76 : data <= 8'b00000000 ;
			15'h00007E77 : data <= 8'b00000000 ;
			15'h00007E78 : data <= 8'b00000000 ;
			15'h00007E79 : data <= 8'b00000000 ;
			15'h00007E7A : data <= 8'b00000000 ;
			15'h00007E7B : data <= 8'b00000000 ;
			15'h00007E7C : data <= 8'b00000000 ;
			15'h00007E7D : data <= 8'b00000000 ;
			15'h00007E7E : data <= 8'b00000000 ;
			15'h00007E7F : data <= 8'b00000000 ;
			15'h00007E80 : data <= 8'b00000000 ;
			15'h00007E81 : data <= 8'b00000000 ;
			15'h00007E82 : data <= 8'b00000000 ;
			15'h00007E83 : data <= 8'b00000000 ;
			15'h00007E84 : data <= 8'b00000000 ;
			15'h00007E85 : data <= 8'b00000000 ;
			15'h00007E86 : data <= 8'b00000000 ;
			15'h00007E87 : data <= 8'b00000000 ;
			15'h00007E88 : data <= 8'b00000000 ;
			15'h00007E89 : data <= 8'b00000000 ;
			15'h00007E8A : data <= 8'b00000000 ;
			15'h00007E8B : data <= 8'b00000000 ;
			15'h00007E8C : data <= 8'b00000000 ;
			15'h00007E8D : data <= 8'b00000000 ;
			15'h00007E8E : data <= 8'b00000000 ;
			15'h00007E8F : data <= 8'b00000000 ;
			15'h00007E90 : data <= 8'b00000000 ;
			15'h00007E91 : data <= 8'b00000000 ;
			15'h00007E92 : data <= 8'b00000000 ;
			15'h00007E93 : data <= 8'b00000000 ;
			15'h00007E94 : data <= 8'b00000000 ;
			15'h00007E95 : data <= 8'b00000000 ;
			15'h00007E96 : data <= 8'b00000000 ;
			15'h00007E97 : data <= 8'b00000000 ;
			15'h00007E98 : data <= 8'b00000000 ;
			15'h00007E99 : data <= 8'b00000000 ;
			15'h00007E9A : data <= 8'b00000000 ;
			15'h00007E9B : data <= 8'b00000000 ;
			15'h00007E9C : data <= 8'b00000000 ;
			15'h00007E9D : data <= 8'b00000000 ;
			15'h00007E9E : data <= 8'b00000000 ;
			15'h00007E9F : data <= 8'b00000000 ;
			15'h00007EA0 : data <= 8'b00000000 ;
			15'h00007EA1 : data <= 8'b00000000 ;
			15'h00007EA2 : data <= 8'b00000000 ;
			15'h00007EA3 : data <= 8'b00000000 ;
			15'h00007EA4 : data <= 8'b00000000 ;
			15'h00007EA5 : data <= 8'b00000000 ;
			15'h00007EA6 : data <= 8'b00000000 ;
			15'h00007EA7 : data <= 8'b00000000 ;
			15'h00007EA8 : data <= 8'b00000000 ;
			15'h00007EA9 : data <= 8'b00000000 ;
			15'h00007EAA : data <= 8'b00000000 ;
			15'h00007EAB : data <= 8'b00000000 ;
			15'h00007EAC : data <= 8'b00000000 ;
			15'h00007EAD : data <= 8'b00000000 ;
			15'h00007EAE : data <= 8'b00000000 ;
			15'h00007EAF : data <= 8'b00000000 ;
			15'h00007EB0 : data <= 8'b00000000 ;
			15'h00007EB1 : data <= 8'b00000000 ;
			15'h00007EB2 : data <= 8'b00000000 ;
			15'h00007EB3 : data <= 8'b00000000 ;
			15'h00007EB4 : data <= 8'b00000000 ;
			15'h00007EB5 : data <= 8'b00000000 ;
			15'h00007EB6 : data <= 8'b00000000 ;
			15'h00007EB7 : data <= 8'b00000000 ;
			15'h00007EB8 : data <= 8'b00000000 ;
			15'h00007EB9 : data <= 8'b00000000 ;
			15'h00007EBA : data <= 8'b00000000 ;
			15'h00007EBB : data <= 8'b00000000 ;
			15'h00007EBC : data <= 8'b00000000 ;
			15'h00007EBD : data <= 8'b00000000 ;
			15'h00007EBE : data <= 8'b00000000 ;
			15'h00007EBF : data <= 8'b00000000 ;
			15'h00007EC0 : data <= 8'b00000000 ;
			15'h00007EC1 : data <= 8'b00000000 ;
			15'h00007EC2 : data <= 8'b00000000 ;
			15'h00007EC3 : data <= 8'b00000000 ;
			15'h00007EC4 : data <= 8'b00000000 ;
			15'h00007EC5 : data <= 8'b00000000 ;
			15'h00007EC6 : data <= 8'b00000000 ;
			15'h00007EC7 : data <= 8'b00000000 ;
			15'h00007EC8 : data <= 8'b00000000 ;
			15'h00007EC9 : data <= 8'b00000000 ;
			15'h00007ECA : data <= 8'b00000000 ;
			15'h00007ECB : data <= 8'b00000000 ;
			15'h00007ECC : data <= 8'b00000000 ;
			15'h00007ECD : data <= 8'b00000000 ;
			15'h00007ECE : data <= 8'b00000000 ;
			15'h00007ECF : data <= 8'b00000000 ;
			15'h00007ED0 : data <= 8'b00000000 ;
			15'h00007ED1 : data <= 8'b00000000 ;
			15'h00007ED2 : data <= 8'b00000000 ;
			15'h00007ED3 : data <= 8'b00000000 ;
			15'h00007ED4 : data <= 8'b00000000 ;
			15'h00007ED5 : data <= 8'b00000000 ;
			15'h00007ED6 : data <= 8'b00000000 ;
			15'h00007ED7 : data <= 8'b00000000 ;
			15'h00007ED8 : data <= 8'b00000000 ;
			15'h00007ED9 : data <= 8'b00000000 ;
			15'h00007EDA : data <= 8'b00000000 ;
			15'h00007EDB : data <= 8'b00000000 ;
			15'h00007EDC : data <= 8'b00000000 ;
			15'h00007EDD : data <= 8'b00000000 ;
			15'h00007EDE : data <= 8'b00000000 ;
			15'h00007EDF : data <= 8'b00000000 ;
			15'h00007EE0 : data <= 8'b00000000 ;
			15'h00007EE1 : data <= 8'b00000000 ;
			15'h00007EE2 : data <= 8'b00000000 ;
			15'h00007EE3 : data <= 8'b00000000 ;
			15'h00007EE4 : data <= 8'b00000000 ;
			15'h00007EE5 : data <= 8'b00000000 ;
			15'h00007EE6 : data <= 8'b00000000 ;
			15'h00007EE7 : data <= 8'b00000000 ;
			15'h00007EE8 : data <= 8'b00000000 ;
			15'h00007EE9 : data <= 8'b00000000 ;
			15'h00007EEA : data <= 8'b00000000 ;
			15'h00007EEB : data <= 8'b00000000 ;
			15'h00007EEC : data <= 8'b00000000 ;
			15'h00007EED : data <= 8'b00000000 ;
			15'h00007EEE : data <= 8'b00000000 ;
			15'h00007EEF : data <= 8'b00000000 ;
			15'h00007EF0 : data <= 8'b00000000 ;
			15'h00007EF1 : data <= 8'b00000000 ;
			15'h00007EF2 : data <= 8'b00000000 ;
			15'h00007EF3 : data <= 8'b00000000 ;
			15'h00007EF4 : data <= 8'b00000000 ;
			15'h00007EF5 : data <= 8'b00000000 ;
			15'h00007EF6 : data <= 8'b00000000 ;
			15'h00007EF7 : data <= 8'b00000000 ;
			15'h00007EF8 : data <= 8'b00000000 ;
			15'h00007EF9 : data <= 8'b00000000 ;
			15'h00007EFA : data <= 8'b00000000 ;
			15'h00007EFB : data <= 8'b00000000 ;
			15'h00007EFC : data <= 8'b00000000 ;
			15'h00007EFD : data <= 8'b00000000 ;
			15'h00007EFE : data <= 8'b00000000 ;
			15'h00007EFF : data <= 8'b00000000 ;
			15'h00007F00 : data <= 8'b00000000 ;
			15'h00007F01 : data <= 8'b00000000 ;
			15'h00007F02 : data <= 8'b00000000 ;
			15'h00007F03 : data <= 8'b00000000 ;
			15'h00007F04 : data <= 8'b00000000 ;
			15'h00007F05 : data <= 8'b00000000 ;
			15'h00007F06 : data <= 8'b00000000 ;
			15'h00007F07 : data <= 8'b00000000 ;
			15'h00007F08 : data <= 8'b00000000 ;
			15'h00007F09 : data <= 8'b00000000 ;
			15'h00007F0A : data <= 8'b00000000 ;
			15'h00007F0B : data <= 8'b00000000 ;
			15'h00007F0C : data <= 8'b00000000 ;
			15'h00007F0D : data <= 8'b00000000 ;
			15'h00007F0E : data <= 8'b00000000 ;
			15'h00007F0F : data <= 8'b00000000 ;
			15'h00007F10 : data <= 8'b00000000 ;
			15'h00007F11 : data <= 8'b00000000 ;
			15'h00007F12 : data <= 8'b00000000 ;
			15'h00007F13 : data <= 8'b00000000 ;
			15'h00007F14 : data <= 8'b00000000 ;
			15'h00007F15 : data <= 8'b00000000 ;
			15'h00007F16 : data <= 8'b00000000 ;
			15'h00007F17 : data <= 8'b00000000 ;
			15'h00007F18 : data <= 8'b00000000 ;
			15'h00007F19 : data <= 8'b00000000 ;
			15'h00007F1A : data <= 8'b00000000 ;
			15'h00007F1B : data <= 8'b00000000 ;
			15'h00007F1C : data <= 8'b00000000 ;
			15'h00007F1D : data <= 8'b00000000 ;
			15'h00007F1E : data <= 8'b00000000 ;
			15'h00007F1F : data <= 8'b00000000 ;
			15'h00007F20 : data <= 8'b00000000 ;
			15'h00007F21 : data <= 8'b00000000 ;
			15'h00007F22 : data <= 8'b00000000 ;
			15'h00007F23 : data <= 8'b00000000 ;
			15'h00007F24 : data <= 8'b00000000 ;
			15'h00007F25 : data <= 8'b00000000 ;
			15'h00007F26 : data <= 8'b00000000 ;
			15'h00007F27 : data <= 8'b00000000 ;
			15'h00007F28 : data <= 8'b00000000 ;
			15'h00007F29 : data <= 8'b00000000 ;
			15'h00007F2A : data <= 8'b00000000 ;
			15'h00007F2B : data <= 8'b00000000 ;
			15'h00007F2C : data <= 8'b00000000 ;
			15'h00007F2D : data <= 8'b00000000 ;
			15'h00007F2E : data <= 8'b00000000 ;
			15'h00007F2F : data <= 8'b00000000 ;
			15'h00007F30 : data <= 8'b00000000 ;
			15'h00007F31 : data <= 8'b00000000 ;
			15'h00007F32 : data <= 8'b00000000 ;
			15'h00007F33 : data <= 8'b00000000 ;
			15'h00007F34 : data <= 8'b00000000 ;
			15'h00007F35 : data <= 8'b00000000 ;
			15'h00007F36 : data <= 8'b00000000 ;
			15'h00007F37 : data <= 8'b00000000 ;
			15'h00007F38 : data <= 8'b00000000 ;
			15'h00007F39 : data <= 8'b00000000 ;
			15'h00007F3A : data <= 8'b00000000 ;
			15'h00007F3B : data <= 8'b00000000 ;
			15'h00007F3C : data <= 8'b00000000 ;
			15'h00007F3D : data <= 8'b00000000 ;
			15'h00007F3E : data <= 8'b00000000 ;
			15'h00007F3F : data <= 8'b00000000 ;
			15'h00007F40 : data <= 8'b00000000 ;
			15'h00007F41 : data <= 8'b00000000 ;
			15'h00007F42 : data <= 8'b00000000 ;
			15'h00007F43 : data <= 8'b00000000 ;
			15'h00007F44 : data <= 8'b00000000 ;
			15'h00007F45 : data <= 8'b00000000 ;
			15'h00007F46 : data <= 8'b00000000 ;
			15'h00007F47 : data <= 8'b00000000 ;
			15'h00007F48 : data <= 8'b00000000 ;
			15'h00007F49 : data <= 8'b00000000 ;
			15'h00007F4A : data <= 8'b00000000 ;
			15'h00007F4B : data <= 8'b00000000 ;
			15'h00007F4C : data <= 8'b00000000 ;
			15'h00007F4D : data <= 8'b00000000 ;
			15'h00007F4E : data <= 8'b00000000 ;
			15'h00007F4F : data <= 8'b00000000 ;
			15'h00007F50 : data <= 8'b00000000 ;
			15'h00007F51 : data <= 8'b00000000 ;
			15'h00007F52 : data <= 8'b00000000 ;
			15'h00007F53 : data <= 8'b00000000 ;
			15'h00007F54 : data <= 8'b00000000 ;
			15'h00007F55 : data <= 8'b00000000 ;
			15'h00007F56 : data <= 8'b00000000 ;
			15'h00007F57 : data <= 8'b00000000 ;
			15'h00007F58 : data <= 8'b00000000 ;
			15'h00007F59 : data <= 8'b00000000 ;
			15'h00007F5A : data <= 8'b00000000 ;
			15'h00007F5B : data <= 8'b00000000 ;
			15'h00007F5C : data <= 8'b00000000 ;
			15'h00007F5D : data <= 8'b00000000 ;
			15'h00007F5E : data <= 8'b00000000 ;
			15'h00007F5F : data <= 8'b00000000 ;
			15'h00007F60 : data <= 8'b00000000 ;
			15'h00007F61 : data <= 8'b00000000 ;
			15'h00007F62 : data <= 8'b00000000 ;
			15'h00007F63 : data <= 8'b00000000 ;
			15'h00007F64 : data <= 8'b00000000 ;
			15'h00007F65 : data <= 8'b00000000 ;
			15'h00007F66 : data <= 8'b00000000 ;
			15'h00007F67 : data <= 8'b00000000 ;
			15'h00007F68 : data <= 8'b00000000 ;
			15'h00007F69 : data <= 8'b00000000 ;
			15'h00007F6A : data <= 8'b00000000 ;
			15'h00007F6B : data <= 8'b00000000 ;
			15'h00007F6C : data <= 8'b00000000 ;
			15'h00007F6D : data <= 8'b00000000 ;
			15'h00007F6E : data <= 8'b00000000 ;
			15'h00007F6F : data <= 8'b00000000 ;
			15'h00007F70 : data <= 8'b00000000 ;
			15'h00007F71 : data <= 8'b00000000 ;
			15'h00007F72 : data <= 8'b00000000 ;
			15'h00007F73 : data <= 8'b00000000 ;
			15'h00007F74 : data <= 8'b00000000 ;
			15'h00007F75 : data <= 8'b00000000 ;
			15'h00007F76 : data <= 8'b00000000 ;
			15'h00007F77 : data <= 8'b00000000 ;
			15'h00007F78 : data <= 8'b00000000 ;
			15'h00007F79 : data <= 8'b00000000 ;
			15'h00007F7A : data <= 8'b00000000 ;
			15'h00007F7B : data <= 8'b00000000 ;
			15'h00007F7C : data <= 8'b00000000 ;
			15'h00007F7D : data <= 8'b00000000 ;
			15'h00007F7E : data <= 8'b00000000 ;
			15'h00007F7F : data <= 8'b00000000 ;
			15'h00007F80 : data <= 8'b00000000 ;
			15'h00007F81 : data <= 8'b00000000 ;
			15'h00007F82 : data <= 8'b00000000 ;
			15'h00007F83 : data <= 8'b00000000 ;
			15'h00007F84 : data <= 8'b00000000 ;
			15'h00007F85 : data <= 8'b00000000 ;
			15'h00007F86 : data <= 8'b00000000 ;
			15'h00007F87 : data <= 8'b00000000 ;
			15'h00007F88 : data <= 8'b00000000 ;
			15'h00007F89 : data <= 8'b00000000 ;
			15'h00007F8A : data <= 8'b00000000 ;
			15'h00007F8B : data <= 8'b00000000 ;
			15'h00007F8C : data <= 8'b00000000 ;
			15'h00007F8D : data <= 8'b00000000 ;
			15'h00007F8E : data <= 8'b00000000 ;
			15'h00007F8F : data <= 8'b00000000 ;
			15'h00007F90 : data <= 8'b00000000 ;
			15'h00007F91 : data <= 8'b00000000 ;
			15'h00007F92 : data <= 8'b00000000 ;
			15'h00007F93 : data <= 8'b00000000 ;
			15'h00007F94 : data <= 8'b00000000 ;
			15'h00007F95 : data <= 8'b00000000 ;
			15'h00007F96 : data <= 8'b00000000 ;
			15'h00007F97 : data <= 8'b00000000 ;
			15'h00007F98 : data <= 8'b00000000 ;
			15'h00007F99 : data <= 8'b00000000 ;
			15'h00007F9A : data <= 8'b00000000 ;
			15'h00007F9B : data <= 8'b00000000 ;
			15'h00007F9C : data <= 8'b00000000 ;
			15'h00007F9D : data <= 8'b00000000 ;
			15'h00007F9E : data <= 8'b00000000 ;
			15'h00007F9F : data <= 8'b00000000 ;
			15'h00007FA0 : data <= 8'b00000000 ;
			15'h00007FA1 : data <= 8'b00000000 ;
			15'h00007FA2 : data <= 8'b00000000 ;
			15'h00007FA3 : data <= 8'b00000000 ;
			15'h00007FA4 : data <= 8'b00000000 ;
			15'h00007FA5 : data <= 8'b00000000 ;
			15'h00007FA6 : data <= 8'b00000000 ;
			15'h00007FA7 : data <= 8'b00000000 ;
			15'h00007FA8 : data <= 8'b00000000 ;
			15'h00007FA9 : data <= 8'b00000000 ;
			15'h00007FAA : data <= 8'b00000000 ;
			15'h00007FAB : data <= 8'b00000000 ;
			15'h00007FAC : data <= 8'b00000000 ;
			15'h00007FAD : data <= 8'b00000000 ;
			15'h00007FAE : data <= 8'b00000000 ;
			15'h00007FAF : data <= 8'b00000000 ;
			15'h00007FB0 : data <= 8'b00000000 ;
			15'h00007FB1 : data <= 8'b00000000 ;
			15'h00007FB2 : data <= 8'b00000000 ;
			15'h00007FB3 : data <= 8'b00000000 ;
			15'h00007FB4 : data <= 8'b00000000 ;
			15'h00007FB5 : data <= 8'b00000000 ;
			15'h00007FB6 : data <= 8'b00000000 ;
			15'h00007FB7 : data <= 8'b00000000 ;
			15'h00007FB8 : data <= 8'b00000000 ;
			15'h00007FB9 : data <= 8'b00000000 ;
			15'h00007FBA : data <= 8'b00000000 ;
			15'h00007FBB : data <= 8'b00000000 ;
			15'h00007FBC : data <= 8'b00000000 ;
			15'h00007FBD : data <= 8'b00000000 ;
			15'h00007FBE : data <= 8'b00000000 ;
			15'h00007FBF : data <= 8'b00000000 ;
			15'h00007FC0 : data <= 8'b00000000 ;
			15'h00007FC1 : data <= 8'b00000000 ;
			15'h00007FC2 : data <= 8'b00000000 ;
			15'h00007FC3 : data <= 8'b00000000 ;
			15'h00007FC4 : data <= 8'b00000000 ;
			15'h00007FC5 : data <= 8'b00000000 ;
			15'h00007FC6 : data <= 8'b00000000 ;
			15'h00007FC7 : data <= 8'b00000000 ;
			15'h00007FC8 : data <= 8'b00000000 ;
			15'h00007FC9 : data <= 8'b00000000 ;
			15'h00007FCA : data <= 8'b00000000 ;
			15'h00007FCB : data <= 8'b00000000 ;
			15'h00007FCC : data <= 8'b00000000 ;
			15'h00007FCD : data <= 8'b00000000 ;
			15'h00007FCE : data <= 8'b00000000 ;
			15'h00007FCF : data <= 8'b00000000 ;
			15'h00007FD0 : data <= 8'b00000000 ;
			15'h00007FD1 : data <= 8'b00000000 ;
			15'h00007FD2 : data <= 8'b00000000 ;
			15'h00007FD3 : data <= 8'b00000000 ;
			15'h00007FD4 : data <= 8'b00000000 ;
			15'h00007FD5 : data <= 8'b00000000 ;
			15'h00007FD6 : data <= 8'b00000000 ;
			15'h00007FD7 : data <= 8'b00000000 ;
			15'h00007FD8 : data <= 8'b00000000 ;
			15'h00007FD9 : data <= 8'b00000000 ;
			15'h00007FDA : data <= 8'b00000000 ;
			15'h00007FDB : data <= 8'b00000000 ;
			15'h00007FDC : data <= 8'b00000000 ;
			15'h00007FDD : data <= 8'b00000000 ;
			15'h00007FDE : data <= 8'b00000000 ;
			15'h00007FDF : data <= 8'b00000000 ;
			15'h00007FE0 : data <= 8'b00000000 ;
			15'h00007FE1 : data <= 8'b00000000 ;
			15'h00007FE2 : data <= 8'b00000000 ;
			15'h00007FE3 : data <= 8'b00000000 ;
			15'h00007FE4 : data <= 8'b00000000 ;
			15'h00007FE5 : data <= 8'b00000000 ;
			15'h00007FE6 : data <= 8'b00000000 ;
			15'h00007FE7 : data <= 8'b00000000 ;
			15'h00007FE8 : data <= 8'b00000000 ;
			15'h00007FE9 : data <= 8'b00000000 ;
			15'h00007FEA : data <= 8'b00000000 ;
			15'h00007FEB : data <= 8'b00000000 ;
			15'h00007FEC : data <= 8'b00000000 ;
			15'h00007FED : data <= 8'b00000000 ;
			15'h00007FEE : data <= 8'b00000000 ;
			15'h00007FEF : data <= 8'b00000000 ;
			15'h00007FF0 : data <= 8'b00000000 ;
			15'h00007FF1 : data <= 8'b00000000 ;
			15'h00007FF2 : data <= 8'b00000000 ;
			15'h00007FF3 : data <= 8'b00000000 ;
			15'h00007FF4 : data <= 8'b00000000 ;
			15'h00007FF5 : data <= 8'b00000000 ;
			15'h00007FF6 : data <= 8'b00000000 ;
			15'h00007FF7 : data <= 8'b00000000 ;
			15'h00007FF8 : data <= 8'b00000000 ;
			15'h00007FF9 : data <= 8'b00000000 ;
			15'h00007FFA : data <= 8'b00000000 ;
			15'h00007FFB : data <= 8'b10000000 ;
			15'h00007FFC : data <= 8'b00000000 ;
			15'h00007FFD : data <= 8'b10000000 ;
			15'h00007FFE : data <= 8'b00000000 ;
			15'h00007FFF : data <= 8'b10000000 ;
		endcase
	end
endmodule