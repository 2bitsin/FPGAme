
module screen0 (clock, addr, data);
	input wire clock;
	input wire[8:0] addr;
	(* romstyle = "M10K" *)
	output bit[7:0] data;
	always @(posedge clock)
	begin
		case(addr)
			9'h00000000 : data <= 8'b00100000 ;
			9'h00000001 : data <= 8'b00100000 ;
			9'h00000002 : data <= 8'b00100000 ;
			9'h00000003 : data <= 8'b00100000 ;
			9'h00000004 : data <= 8'b00100000 ;
			9'h00000005 : data <= 8'b00100000 ;
			9'h00000006 : data <= 8'b00100000 ;
			9'h00000007 : data <= 8'b00100000 ;
			9'h00000008 : data <= 8'b00100000 ;
			9'h00000009 : data <= 8'b00100000 ;
			9'h0000000A : data <= 8'b00100000 ;
			9'h0000000B : data <= 8'b00100000 ;
			9'h0000000C : data <= 8'b00100000 ;
			9'h0000000D : data <= 8'b00100000 ;
			9'h0000000E : data <= 8'b00100000 ;
			9'h0000000F : data <= 8'b00100000 ;
			9'h00000010 : data <= 8'b00100000 ;
			9'h00000011 : data <= 8'b00100000 ;
			9'h00000012 : data <= 8'b00100000 ;
			9'h00000013 : data <= 8'b00100000 ;
			9'h00000014 : data <= 8'b00100000 ;
			9'h00000015 : data <= 8'b00100000 ;
			9'h00000016 : data <= 8'b00100000 ;
			9'h00000017 : data <= 8'b00100000 ;
			9'h00000018 : data <= 8'b00100000 ;
			9'h00000019 : data <= 8'b00100000 ;
			9'h0000001A : data <= 8'b00100000 ;
			9'h0000001B : data <= 8'b00100000 ;
			9'h0000001C : data <= 8'b00100000 ;
			9'h0000001D : data <= 8'b00100000 ;
			9'h0000001E : data <= 8'b00100000 ;
			9'h0000001F : data <= 8'b00100000 ;
			9'h00000020 : data <= 8'b00100000 ;
			9'h00000021 : data <= 8'b00100000 ;
			9'h00000022 : data <= 8'b00100000 ;
			9'h00000023 : data <= 8'b00100000 ;
			9'h00000024 : data <= 8'b00100000 ;
			9'h00000025 : data <= 8'b00100000 ;
			9'h00000026 : data <= 8'b00100000 ;
			9'h00000027 : data <= 8'b00100000 ;
			9'h00000028 : data <= 8'b00100000 ;
			9'h00000029 : data <= 8'b00100000 ;
			9'h0000002A : data <= 8'b00100000 ;
			9'h0000002B : data <= 8'b00100000 ;
			9'h0000002C : data <= 8'b00100000 ;
			9'h0000002D : data <= 8'b00100000 ;
			9'h0000002E : data <= 8'b00100000 ;
			9'h0000002F : data <= 8'b00100000 ;
			9'h00000030 : data <= 8'b00100000 ;
			9'h00000031 : data <= 8'b00100000 ;
			9'h00000032 : data <= 8'b00100000 ;
			9'h00000033 : data <= 8'b00100000 ;
			9'h00000034 : data <= 8'b00100000 ;
			9'h00000035 : data <= 8'b00100000 ;
			9'h00000036 : data <= 8'b00100000 ;
			9'h00000037 : data <= 8'b00100000 ;
			9'h00000038 : data <= 8'b00100000 ;
			9'h00000039 : data <= 8'b00100000 ;
			9'h0000003A : data <= 8'b00100000 ;
			9'h0000003B : data <= 8'b00100000 ;
			9'h0000003C : data <= 8'b00100000 ;
			9'h0000003D : data <= 8'b00100000 ;
			9'h0000003E : data <= 8'b00100000 ;
			9'h0000003F : data <= 8'b00100000 ;
			9'h00000040 : data <= 8'b00100000 ;
			9'h00000041 : data <= 8'b00100000 ;
			9'h00000042 : data <= 8'b00101011 ;
			9'h00000043 : data <= 8'b00101101 ;
			9'h00000044 : data <= 8'b00101101 ;
			9'h00000045 : data <= 8'b00101101 ;
			9'h00000046 : data <= 8'b00101101 ;
			9'h00000047 : data <= 8'b00101101 ;
			9'h00000048 : data <= 8'b00101101 ;
			9'h00000049 : data <= 8'b00101101 ;
			9'h0000004A : data <= 8'b00101101 ;
			9'h0000004B : data <= 8'b00101101 ;
			9'h0000004C : data <= 8'b00101101 ;
			9'h0000004D : data <= 8'b00101101 ;
			9'h0000004E : data <= 8'b00101101 ;
			9'h0000004F : data <= 8'b00101101 ;
			9'h00000050 : data <= 8'b00101101 ;
			9'h00000051 : data <= 8'b00101101 ;
			9'h00000052 : data <= 8'b00101101 ;
			9'h00000053 : data <= 8'b00101101 ;
			9'h00000054 : data <= 8'b00101101 ;
			9'h00000055 : data <= 8'b00101101 ;
			9'h00000056 : data <= 8'b00101101 ;
			9'h00000057 : data <= 8'b00101101 ;
			9'h00000058 : data <= 8'b00101101 ;
			9'h00000059 : data <= 8'b00101101 ;
			9'h0000005A : data <= 8'b00101101 ;
			9'h0000005B : data <= 8'b00101101 ;
			9'h0000005C : data <= 8'b00101011 ;
			9'h0000005D : data <= 8'b00100000 ;
			9'h0000005E : data <= 8'b00100000 ;
			9'h0000005F : data <= 8'b00100000 ;
			9'h00000060 : data <= 8'b00100000 ;
			9'h00000061 : data <= 8'b00100000 ;
			9'h00000062 : data <= 8'b01111100 ;
			9'h00000063 : data <= 8'b00100000 ;
			9'h00000064 : data <= 8'b00100000 ;
			9'h00000065 : data <= 8'b00100000 ;
			9'h00000066 : data <= 8'b00100000 ;
			9'h00000067 : data <= 8'b00100000 ;
			9'h00000068 : data <= 8'b00100000 ;
			9'h00000069 : data <= 8'b00100000 ;
			9'h0000006A : data <= 8'b00100000 ;
			9'h0000006B : data <= 8'b00100000 ;
			9'h0000006C : data <= 8'b00100000 ;
			9'h0000006D : data <= 8'b00100000 ;
			9'h0000006E : data <= 8'b00100000 ;
			9'h0000006F : data <= 8'b00100000 ;
			9'h00000070 : data <= 8'b00100000 ;
			9'h00000071 : data <= 8'b00100000 ;
			9'h00000072 : data <= 8'b00100000 ;
			9'h00000073 : data <= 8'b00100000 ;
			9'h00000074 : data <= 8'b00100000 ;
			9'h00000075 : data <= 8'b00100000 ;
			9'h00000076 : data <= 8'b00100000 ;
			9'h00000077 : data <= 8'b00100000 ;
			9'h00000078 : data <= 8'b00100000 ;
			9'h00000079 : data <= 8'b00100000 ;
			9'h0000007A : data <= 8'b00100000 ;
			9'h0000007B : data <= 8'b00100000 ;
			9'h0000007C : data <= 8'b01111100 ;
			9'h0000007D : data <= 8'b00100000 ;
			9'h0000007E : data <= 8'b00100000 ;
			9'h0000007F : data <= 8'b00100000 ;
			9'h00000080 : data <= 8'b00100000 ;
			9'h00000081 : data <= 8'b00100000 ;
			9'h00000082 : data <= 8'b01111100 ;
			9'h00000083 : data <= 8'b00100000 ;
			9'h00000084 : data <= 8'b00100000 ;
			9'h00000085 : data <= 8'b00100000 ;
			9'h00000086 : data <= 8'b00100000 ;
			9'h00000087 : data <= 8'b00100000 ;
			9'h00000088 : data <= 8'b00100000 ;
			9'h00000089 : data <= 8'b00100000 ;
			9'h0000008A : data <= 8'b01001000 ;
			9'h0000008B : data <= 8'b01000101 ;
			9'h0000008C : data <= 8'b01001100 ;
			9'h0000008D : data <= 8'b01001100 ;
			9'h0000008E : data <= 8'b01001111 ;
			9'h0000008F : data <= 8'b00100000 ;
			9'h00000090 : data <= 8'b01010111 ;
			9'h00000091 : data <= 8'b01001111 ;
			9'h00000092 : data <= 8'b01010010 ;
			9'h00000093 : data <= 8'b01001100 ;
			9'h00000094 : data <= 8'b01000100 ;
			9'h00000095 : data <= 8'b00100001 ;
			9'h00000096 : data <= 8'b00100000 ;
			9'h00000097 : data <= 8'b00100000 ;
			9'h00000098 : data <= 8'b00100000 ;
			9'h00000099 : data <= 8'b00100000 ;
			9'h0000009A : data <= 8'b00100000 ;
			9'h0000009B : data <= 8'b00100000 ;
			9'h0000009C : data <= 8'b01111100 ;
			9'h0000009D : data <= 8'b00100000 ;
			9'h0000009E : data <= 8'b00100000 ;
			9'h0000009F : data <= 8'b00100000 ;
			9'h000000A0 : data <= 8'b00100000 ;
			9'h000000A1 : data <= 8'b00100000 ;
			9'h000000A2 : data <= 8'b01111100 ;
			9'h000000A3 : data <= 8'b00100000 ;
			9'h000000A4 : data <= 8'b00100000 ;
			9'h000000A5 : data <= 8'b00100000 ;
			9'h000000A6 : data <= 8'b00100000 ;
			9'h000000A7 : data <= 8'b00100000 ;
			9'h000000A8 : data <= 8'b00100000 ;
			9'h000000A9 : data <= 8'b00100000 ;
			9'h000000AA : data <= 8'b00100000 ;
			9'h000000AB : data <= 8'b00100000 ;
			9'h000000AC : data <= 8'b00100000 ;
			9'h000000AD : data <= 8'b00100000 ;
			9'h000000AE : data <= 8'b01100001 ;
			9'h000000AF : data <= 8'b01101100 ;
			9'h000000B0 : data <= 8'b01100101 ;
			9'h000000B1 : data <= 8'b01111000 ;
			9'h000000B2 : data <= 8'b00100000 ;
			9'h000000B3 : data <= 8'b01101000 ;
			9'h000000B4 : data <= 8'b01100101 ;
			9'h000000B5 : data <= 8'b01110010 ;
			9'h000000B6 : data <= 8'b01100101 ;
			9'h000000B7 : data <= 8'b00101110 ;
			9'h000000B8 : data <= 8'b00101110 ;
			9'h000000B9 : data <= 8'b00100000 ;
			9'h000000BA : data <= 8'b00100000 ;
			9'h000000BB : data <= 8'b00100000 ;
			9'h000000BC : data <= 8'b01111100 ;
			9'h000000BD : data <= 8'b00100000 ;
			9'h000000BE : data <= 8'b00100000 ;
			9'h000000BF : data <= 8'b00100000 ;
			9'h000000C0 : data <= 8'b00100000 ;
			9'h000000C1 : data <= 8'b00100000 ;
			9'h000000C2 : data <= 8'b01111100 ;
			9'h000000C3 : data <= 8'b00100000 ;
			9'h000000C4 : data <= 8'b00100000 ;
			9'h000000C5 : data <= 8'b00100000 ;
			9'h000000C6 : data <= 8'b00100000 ;
			9'h000000C7 : data <= 8'b00100000 ;
			9'h000000C8 : data <= 8'b00100000 ;
			9'h000000C9 : data <= 8'b00100000 ;
			9'h000000CA : data <= 8'b00100000 ;
			9'h000000CB : data <= 8'b00100000 ;
			9'h000000CC : data <= 8'b00100000 ;
			9'h000000CD : data <= 8'b00100000 ;
			9'h000000CE : data <= 8'b00100000 ;
			9'h000000CF : data <= 8'b00100000 ;
			9'h000000D0 : data <= 8'b00100000 ;
			9'h000000D1 : data <= 8'b00100000 ;
			9'h000000D2 : data <= 8'b00100000 ;
			9'h000000D3 : data <= 8'b00100000 ;
			9'h000000D4 : data <= 8'b00100000 ;
			9'h000000D5 : data <= 8'b00100000 ;
			9'h000000D6 : data <= 8'b00100000 ;
			9'h000000D7 : data <= 8'b00100000 ;
			9'h000000D8 : data <= 8'b00100000 ;
			9'h000000D9 : data <= 8'b00100000 ;
			9'h000000DA : data <= 8'b00100000 ;
			9'h000000DB : data <= 8'b00100000 ;
			9'h000000DC : data <= 8'b01111100 ;
			9'h000000DD : data <= 8'b00100000 ;
			9'h000000DE : data <= 8'b00100000 ;
			9'h000000DF : data <= 8'b00100000 ;
			9'h000000E0 : data <= 8'b00100000 ;
			9'h000000E1 : data <= 8'b00100000 ;
			9'h000000E2 : data <= 8'b00101011 ;
			9'h000000E3 : data <= 8'b00101101 ;
			9'h000000E4 : data <= 8'b00101101 ;
			9'h000000E5 : data <= 8'b00101101 ;
			9'h000000E6 : data <= 8'b00101101 ;
			9'h000000E7 : data <= 8'b00101101 ;
			9'h000000E8 : data <= 8'b00101101 ;
			9'h000000E9 : data <= 8'b00101101 ;
			9'h000000EA : data <= 8'b00101101 ;
			9'h000000EB : data <= 8'b00101101 ;
			9'h000000EC : data <= 8'b00101101 ;
			9'h000000ED : data <= 8'b00101101 ;
			9'h000000EE : data <= 8'b00101101 ;
			9'h000000EF : data <= 8'b00101101 ;
			9'h000000F0 : data <= 8'b00101101 ;
			9'h000000F1 : data <= 8'b00101101 ;
			9'h000000F2 : data <= 8'b00101101 ;
			9'h000000F3 : data <= 8'b00101101 ;
			9'h000000F4 : data <= 8'b00101101 ;
			9'h000000F5 : data <= 8'b00101101 ;
			9'h000000F6 : data <= 8'b00101101 ;
			9'h000000F7 : data <= 8'b00101101 ;
			9'h000000F8 : data <= 8'b00101101 ;
			9'h000000F9 : data <= 8'b00101101 ;
			9'h000000FA : data <= 8'b00101101 ;
			9'h000000FB : data <= 8'b00101101 ;
			9'h000000FC : data <= 8'b00101011 ;
			9'h000000FD : data <= 8'b00100000 ;
			9'h000000FE : data <= 8'b00100000 ;
			9'h000000FF : data <= 8'b00100000 ;
			9'h00000100 : data <= 8'b00100000 ;
			9'h00000101 : data <= 8'b00100000 ;
			9'h00000102 : data <= 8'b00100000 ;
			9'h00000103 : data <= 8'b00100000 ;
			9'h00000104 : data <= 8'b00100000 ;
			9'h00000105 : data <= 8'b00100000 ;
			9'h00000106 : data <= 8'b00100000 ;
			9'h00000107 : data <= 8'b00100000 ;
			9'h00000108 : data <= 8'b00100000 ;
			9'h00000109 : data <= 8'b00100000 ;
			9'h0000010A : data <= 8'b10110000 ;
			9'h0000010B : data <= 8'b10110000 ;
			9'h0000010C : data <= 8'b10110000 ;
			9'h0000010D : data <= 8'b10110001 ;
			9'h0000010E : data <= 8'b10110001 ;
			9'h0000010F : data <= 8'b10110001 ;
			9'h00000110 : data <= 8'b10110010 ;
			9'h00000111 : data <= 8'b10110010 ;
			9'h00000112 : data <= 8'b10110010 ;
			9'h00000113 : data <= 8'b00100000 ;
			9'h00000114 : data <= 8'b00100000 ;
			9'h00000115 : data <= 8'b00100000 ;
			9'h00000116 : data <= 8'b00100000 ;
			9'h00000117 : data <= 8'b00100000 ;
			9'h00000118 : data <= 8'b00100000 ;
			9'h00000119 : data <= 8'b00100000 ;
			9'h0000011A : data <= 8'b00100000 ;
			9'h0000011B : data <= 8'b00100000 ;
			9'h0000011C : data <= 8'b00100000 ;
			9'h0000011D : data <= 8'b00100000 ;
			9'h0000011E : data <= 8'b00100000 ;
			9'h0000011F : data <= 8'b00100000 ;
			9'h00000120 : data <= 8'b00100000 ;
			9'h00000121 : data <= 8'b00100000 ;
			9'h00000122 : data <= 8'b00100000 ;
			9'h00000123 : data <= 8'b00100000 ;
			9'h00000124 : data <= 8'b00100000 ;
			9'h00000125 : data <= 8'b00100000 ;
			9'h00000126 : data <= 8'b00100000 ;
			9'h00000127 : data <= 8'b00100000 ;
			9'h00000128 : data <= 8'b00100000 ;
			9'h00000129 : data <= 8'b00100000 ;
			9'h0000012A : data <= 8'b00100000 ;
			9'h0000012B : data <= 8'b00100000 ;
			9'h0000012C : data <= 8'b00100000 ;
			9'h0000012D : data <= 8'b00100000 ;
			9'h0000012E : data <= 8'b00100000 ;
			9'h0000012F : data <= 8'b00100000 ;
			9'h00000130 : data <= 8'b00100000 ;
			9'h00000131 : data <= 8'b00100000 ;
			9'h00000132 : data <= 8'b00100000 ;
			9'h00000133 : data <= 8'b00100000 ;
			9'h00000134 : data <= 8'b00100000 ;
			9'h00000135 : data <= 8'b00100000 ;
			9'h00000136 : data <= 8'b00100000 ;
			9'h00000137 : data <= 8'b00100000 ;
			9'h00000138 : data <= 8'b00100000 ;
			9'h00000139 : data <= 8'b00100000 ;
			9'h0000013A : data <= 8'b00100000 ;
			9'h0000013B : data <= 8'b00100000 ;
			9'h0000013C : data <= 8'b00100000 ;
			9'h0000013D : data <= 8'b00100000 ;
			9'h0000013E : data <= 8'b00100000 ;
			9'h0000013F : data <= 8'b00100000 ;
			9'h00000140 : data <= 8'b00100000 ;
			9'h00000141 : data <= 8'b00100000 ;
			9'h00000142 : data <= 8'b00100000 ;
			9'h00000143 : data <= 8'b00100000 ;
			9'h00000144 : data <= 8'b00100000 ;
			9'h00000145 : data <= 8'b00100000 ;
			9'h00000146 : data <= 8'b00100000 ;
			9'h00000147 : data <= 8'b00100000 ;
			9'h00000148 : data <= 8'b00100000 ;
			9'h00000149 : data <= 8'b00100000 ;
			9'h0000014A : data <= 8'b00100000 ;
			9'h0000014B : data <= 8'b00100000 ;
			9'h0000014C : data <= 8'b00100000 ;
			9'h0000014D : data <= 8'b00100000 ;
			9'h0000014E : data <= 8'b00100000 ;
			9'h0000014F : data <= 8'b00100000 ;
			9'h00000150 : data <= 8'b00100000 ;
			9'h00000151 : data <= 8'b00100000 ;
			9'h00000152 : data <= 8'b00100000 ;
			9'h00000153 : data <= 8'b00100000 ;
			9'h00000154 : data <= 8'b00100000 ;
			9'h00000155 : data <= 8'b00100000 ;
			9'h00000156 : data <= 8'b00100000 ;
			9'h00000157 : data <= 8'b00100000 ;
			9'h00000158 : data <= 8'b00100000 ;
			9'h00000159 : data <= 8'b00100000 ;
			9'h0000015A : data <= 8'b00100000 ;
			9'h0000015B : data <= 8'b00100000 ;
			9'h0000015C : data <= 8'b00100000 ;
			9'h0000015D : data <= 8'b00100000 ;
			9'h0000015E : data <= 8'b00100000 ;
			9'h0000015F : data <= 8'b00100000 ;
			9'h00000160 : data <= 8'b00100000 ;
			9'h00000161 : data <= 8'b00100000 ;
			9'h00000162 : data <= 8'b00100000 ;
			9'h00000163 : data <= 8'b00100000 ;
			9'h00000164 : data <= 8'b00100000 ;
			9'h00000165 : data <= 8'b00100000 ;
			9'h00000166 : data <= 8'b00100000 ;
			9'h00000167 : data <= 8'b00100000 ;
			9'h00000168 : data <= 8'b00100000 ;
			9'h00000169 : data <= 8'b00100000 ;
			9'h0000016A : data <= 8'b00100000 ;
			9'h0000016B : data <= 8'b00100000 ;
			9'h0000016C : data <= 8'b00100000 ;
			9'h0000016D : data <= 8'b00100000 ;
			9'h0000016E : data <= 8'b00100000 ;
			9'h0000016F : data <= 8'b00100000 ;
			9'h00000170 : data <= 8'b00100000 ;
			9'h00000171 : data <= 8'b00100000 ;
			9'h00000172 : data <= 8'b00100000 ;
			9'h00000173 : data <= 8'b00100000 ;
			9'h00000174 : data <= 8'b00100000 ;
			9'h00000175 : data <= 8'b00100000 ;
			9'h00000176 : data <= 8'b00100000 ;
			9'h00000177 : data <= 8'b00100000 ;
			9'h00000178 : data <= 8'b00100000 ;
			9'h00000179 : data <= 8'b00100000 ;
			9'h0000017A : data <= 8'b00100000 ;
			9'h0000017B : data <= 8'b00100000 ;
			9'h0000017C : data <= 8'b00100000 ;
			9'h0000017D : data <= 8'b00100000 ;
			9'h0000017E : data <= 8'b00100000 ;
			9'h0000017F : data <= 8'b00100000 ;
			9'h00000180 : data <= 8'b00100000 ;
			9'h00000181 : data <= 8'b00100000 ;
			9'h00000182 : data <= 8'b00100000 ;
			9'h00000183 : data <= 8'b00100000 ;
			9'h00000184 : data <= 8'b00100000 ;
			9'h00000185 : data <= 8'b00100000 ;
			9'h00000186 : data <= 8'b00100000 ;
			9'h00000187 : data <= 8'b00100000 ;
			9'h00000188 : data <= 8'b00100000 ;
			9'h00000189 : data <= 8'b00100000 ;
			9'h0000018A : data <= 8'b00100000 ;
			9'h0000018B : data <= 8'b00100000 ;
			9'h0000018C : data <= 8'b00100000 ;
			9'h0000018D : data <= 8'b00100000 ;
			9'h0000018E : data <= 8'b00100000 ;
			9'h0000018F : data <= 8'b00100000 ;
			9'h00000190 : data <= 8'b00100000 ;
			9'h00000191 : data <= 8'b00100000 ;
			9'h00000192 : data <= 8'b00100000 ;
			9'h00000193 : data <= 8'b00100000 ;
			9'h00000194 : data <= 8'b00100000 ;
			9'h00000195 : data <= 8'b00100000 ;
			9'h00000196 : data <= 8'b00100000 ;
			9'h00000197 : data <= 8'b00100000 ;
			9'h00000198 : data <= 8'b00100000 ;
			9'h00000199 : data <= 8'b00100000 ;
			9'h0000019A : data <= 8'b00100000 ;
			9'h0000019B : data <= 8'b00100000 ;
			9'h0000019C : data <= 8'b00100000 ;
			9'h0000019D : data <= 8'b00100000 ;
			9'h0000019E : data <= 8'b00100000 ;
			9'h0000019F : data <= 8'b00100000 ;
			9'h000001A0 : data <= 8'b00100000 ;
			9'h000001A1 : data <= 8'b00100000 ;
			9'h000001A2 : data <= 8'b00100000 ;
			9'h000001A3 : data <= 8'b00100000 ;
			9'h000001A4 : data <= 8'b00100000 ;
			9'h000001A5 : data <= 8'b00100000 ;
			9'h000001A6 : data <= 8'b00100000 ;
			9'h000001A7 : data <= 8'b00100000 ;
			9'h000001A8 : data <= 8'b00100000 ;
			9'h000001A9 : data <= 8'b00100000 ;
			9'h000001AA : data <= 8'b00100000 ;
			9'h000001AB : data <= 8'b00100000 ;
			9'h000001AC : data <= 8'b00100000 ;
			9'h000001AD : data <= 8'b00100000 ;
			9'h000001AE : data <= 8'b00100000 ;
			9'h000001AF : data <= 8'b00100000 ;
			9'h000001B0 : data <= 8'b00100000 ;
			9'h000001B1 : data <= 8'b00100000 ;
			9'h000001B2 : data <= 8'b00100000 ;
			9'h000001B3 : data <= 8'b00100000 ;
			9'h000001B4 : data <= 8'b00100000 ;
			9'h000001B5 : data <= 8'b00100000 ;
			9'h000001B6 : data <= 8'b00100000 ;
			9'h000001B7 : data <= 8'b00100000 ;
			9'h000001B8 : data <= 8'b00100000 ;
			9'h000001B9 : data <= 8'b00100000 ;
			9'h000001BA : data <= 8'b00100000 ;
			9'h000001BB : data <= 8'b00100000 ;
			9'h000001BC : data <= 8'b00100000 ;
			9'h000001BD : data <= 8'b00100000 ;
			9'h000001BE : data <= 8'b00100000 ;
			9'h000001BF : data <= 8'b00100000 ;
			9'h000001C0 : data <= 8'b00100000 ;
			9'h000001C1 : data <= 8'b00100000 ;
			9'h000001C2 : data <= 8'b00100000 ;
			9'h000001C3 : data <= 8'b00100000 ;
			9'h000001C4 : data <= 8'b00100000 ;
			9'h000001C5 : data <= 8'b00100000 ;
			9'h000001C6 : data <= 8'b00100000 ;
			9'h000001C7 : data <= 8'b00100000 ;
			9'h000001C8 : data <= 8'b00100000 ;
			9'h000001C9 : data <= 8'b00100000 ;
			9'h000001CA : data <= 8'b00100000 ;
			9'h000001CB : data <= 8'b00100000 ;
			9'h000001CC : data <= 8'b00100000 ;
			9'h000001CD : data <= 8'b00100000 ;
			9'h000001CE : data <= 8'b00100000 ;
			9'h000001CF : data <= 8'b00100000 ;
			9'h000001D0 : data <= 8'b00100000 ;
			9'h000001D1 : data <= 8'b00100000 ;
			9'h000001D2 : data <= 8'b00100000 ;
			9'h000001D3 : data <= 8'b00100000 ;
			9'h000001D4 : data <= 8'b00100000 ;
			9'h000001D5 : data <= 8'b00100000 ;
			9'h000001D6 : data <= 8'b00100000 ;
			9'h000001D7 : data <= 8'b00100000 ;
			9'h000001D8 : data <= 8'b00100000 ;
			9'h000001D9 : data <= 8'b00100000 ;
			9'h000001DA : data <= 8'b00100000 ;
			9'h000001DB : data <= 8'b00100000 ;
			9'h000001DC : data <= 8'b00100000 ;
			9'h000001DD : data <= 8'b00100000 ;
			9'h000001DE : data <= 8'b00100000 ;
			9'h000001DF : data <= 8'b00100000 ;
			9'h000001E0 : data <= 8'b00100000 ;
			9'h000001E1 : data <= 8'b00100000 ;
			9'h000001E2 : data <= 8'b00100000 ;
			9'h000001E3 : data <= 8'b00100000 ;
			9'h000001E4 : data <= 8'b00100000 ;
			9'h000001E5 : data <= 8'b00100000 ;
			9'h000001E6 : data <= 8'b00100000 ;
			9'h000001E7 : data <= 8'b00100000 ;
			9'h000001E8 : data <= 8'b00100000 ;
			9'h000001E9 : data <= 8'b00100000 ;
			9'h000001EA : data <= 8'b00100000 ;
			9'h000001EB : data <= 8'b00100000 ;
			9'h000001EC : data <= 8'b00100000 ;
			9'h000001ED : data <= 8'b00100000 ;
			9'h000001EE : data <= 8'b00100000 ;
			9'h000001EF : data <= 8'b00100000 ;
			9'h000001F0 : data <= 8'b00100000 ;
			9'h000001F1 : data <= 8'b00100000 ;
			9'h000001F2 : data <= 8'b00100000 ;
			9'h000001F3 : data <= 8'b00100000 ;
			9'h000001F4 : data <= 8'b00100000 ;
			9'h000001F5 : data <= 8'b00100000 ;
			9'h000001F6 : data <= 8'b00100000 ;
			9'h000001F7 : data <= 8'b00100000 ;
			9'h000001F8 : data <= 8'b00100000 ;
			9'h000001F9 : data <= 8'b00100000 ;
			9'h000001FA : data <= 8'b00100000 ;
			9'h000001FB : data <= 8'b00100000 ;
			9'h000001FC : data <= 8'b00100000 ;
			9'h000001FD : data <= 8'b00100000 ;
			9'h000001FE : data <= 8'b00100000 ;
			9'h000001FF : data <= 8'b00100000 ;			
		endcase
	end
endmodule